PK   ¬eX�n�  �     cirkitFile.json�][o�:�+�e�*Jy<8�@Ξ�>$�!Kr#�k�����Kʗĺ84�q��Cш��p�qn)ߣM��Z͊���}�6�z��n��D�������&�c��5���M���|w��ͷ�*.֟׫j��*)WsW��JY��ŉ`Y��y�
=c����$x:Ǧl�Ħ+l�Ʀ'�t�MO�陝�<y���r��8��|���\ĥɪXe&�s)M���-ʲ��23n�G@��D-a�A�r�\��'����A�s�<m����]@w��9tw��	��	�c����ܽ�=��'w�t>�J�K�r`�x+�����$�*�)�8S��UUdq&X���{����. :��ڻ^7�v���r.�Kq\{�r��l`�6b_;��]��1�K�\{�c\�v��%*!v���|=�����t�s��.���C.����\{7Ŀ|�(��r|=A�Aq�,X?��e��y{�(����@Y�]�wM�ZB��I�gH|���3��N2��]����]���u��:�gDs�4�3,�N��ө�)��㳏b�\o�g��Y���� �"I�(.��KB�ŐpII�d��b�IS!�#/z9|9~9�y������#lh �i0�i@�3��G1�J!l�(6��`ʖM^AGSРXРX��aA�bA�bѢ8ӌ�����<��=ZV�#
Fl,,	z`0t(���4���TU��H{��Z7�DjذU�i$"b��B ���	��Hd�cà�-�D)��	�*�D��hSqb��xXՕH&2�Mŉ�f
aY"�Ȍ7'��aHd"��c	QX��|4�[�=���b�� �E��9�ou�|Z�[�$Ю~-T�-[�������칐�m�B�����K���s$\$	E�E�pIH�.)	��uD�A/��/��/�0�A0��0��0�1�A��A� ��4(4(4(4(4(4(4(#(+$0�T��XXVH$�h�t�I$9�a�D�F�|X!�D��VH$�h��I$1ja�D�F�cX!�D""S˩��:��H#��&��c�}`!�F&2�Mŉ����D���7'6�φ�ޅD�˫9�w!��j�]HĹ��xq./�돉���f׏8�˯���K�����e^T�^�֛��D7�Toa��~B�FFX�3�)%h��A�K��	��ᦧ覧�����KO���cK�����q��1�ȦKl�
]9�ɠMG݋D�>��K�T�v�66�/BK���t���ub�7�����A����l��|U��Vη�:���oh��$h���O
�d���0��U��@� ����;�g=��5���LI�z2��Ӧ7�	��D�����I��"��
�Y��M�p@�Y$� �-\Y�"��@xF�0��'* ���«��������~O���f}�}�XD�짺D;�g`�52_��%8_��58?�p~
�w� ��g�+�7UCxD�QDr��d�(��$z�(H9�R�´햆�����%��?���}	E�@Q,P�*P�
�m�tgS�e��B� �����i��GaM����-
5p(	�� 
%_�a=ӠP���6
�`��.�I��	��2��}aӠP�4���!�[5�V������hTӌ�`�~`�3*��y�{�Q9�n?a	�l	��{��$���B��.�sA@@��9�����~ F*�)}�N��ԥ+�Y�[W�����a���s�9�uq���ܳM�P�����;R�h�#n��#��s7����h�:�w�f7C���n�p3v�����B���>�������=����E���C��1rr����AA?��'�nؾIC���XX���o�ѯ�CJ�c��
��C�<��&�_�G���ճ�nܫ=�|^-������_U�7'j���C�?$�C�?$�C�?��C�?��C�?d�C�y�|���؇z�Xϖ��i�צ����3_n��̲i��G�4�ӓ�̞.����-���7�����������4u�����n�?�{����4M�T-o3�BNS��2斱Ի�*U�Y�`E�s#�/X�r���y���ێ� ���$�Q���#��h�7��懶�*-�zS,��oe�z"$���&"�e9�����u�4(��_���uƧB&L��u#�*U���|��S#9g"�+k]�if��s�'Sa����u��S��d纱�s��\�V�D�������t*���AJ��U�d?�LN��.�sg��(��wh�����א�f�p���۝�g�KͳsTn�Չ:ǫ�f�g��Ia�� � �ݯD�v����Tv��T��Rٽ�<I�qo����J�l��d��n��:�ь��}O���?�J��H��Y*	�H��g��Pi��p�sp1���=\,��d��Q�O�|h��z}��ʩ���U�*{~�D�v�5-i�w.�A�V��iib{X�1�"fs��e9/yQsST�It�W��5H�j��L���$�� ���Tk�u��:܏�q��Nm�yĴsR���kiK���h��#ֈ�cX�	o�mXwD���^��[���iU��m�~�#�VM�`���[m�D��{TR粿�e��k�T��MO���#��^4Y��~�L�v����y�P�����M�4����/�vo�8���.j�F��n�<��&w���M�^�+�!$�l�U�r�ۥ�g�j���t��i��!_)g���t�>��U�>oZ^����"���x�>4�z�q��ܺ�� ;�(3�^�,�`�RYK@��G�����E?,�~�x���拔Kd�*6� �L_^��R�S<�����Ǎj��Wb@%t�G_O	�����y�O��~v����~9�x���b˓RX�a(@5bS�!�������>M(C�+z2C�'G&7W�Tv��r��K�d�ꗃ�_���p�ud	�#J�E�Q������G5B���E�E^(�(� (���2�T�:����~9�x>l�&R�#F�F@����C5�˰�%T��V�GC�%� ů�lIb@�l��d89�Rf���y����ׇ�ߣ�k"��I	
'5#D �I}�I��Ɯ��sF�@�N�_)b�i��)����a�sJ��p<sx��\B�iS�*~*�D
�M	Jצ�k-<�^>��)=�1��?�FN�+ƽ�(Aao(�
���z�I�ps={������a��\xlo�j,9�z�K�F�{d^/�.�țjS��mt�гm��[�䫧|���ӻ���u����PK   �eX��D>  ?>  /   images/3d2da6db-3dc1-43d2-90bb-751371ef683b.png?>���PNG

   IHDR   d   �   (�-F   	pHYs  ��  �����   tEXtSoftware www.inkscape.org��<  =�IDATx��}x�u�?3��ŢW�;ER%QT�:-Q�r��{�{lŶ�����;Q���ʲ;J,ٲ��%J�D�)���lߙy�3�X� � Rrx���3;3���Ϲ�����6Y�H���K��W�৯� �� M�m[�/���%���q�?�o\W�eeAܳw �n��-�Ć�����߄������x�=�]�q�N�<,|�
�ǎ^ܱ��H���P���ڃ�T��>�����R���`wW#㺤.���_�i�}^U���룿oD����?Z�C}1lk���4>�6���˱q� ��B'.^P�Ｅ^��?f�}�(j�eM9n{�	[[G��˪q��R�b{݁SʲqaM>��H��6 a����m�l.JJ'W/*�W���gj�ֶ(���Q�0zQ��T:GS��LbOw����͈���{����rܷߺ�߹��!�:2��܃=�yZ���,Ë�a������\���X+�m
��7�"����>�'���a���c�o�`4��ҧ&��2�no.�y]5�ws=��a���](Т��>��>75���o���\��է���������a��"L��B �[F��&�z��De�$�f`���\|��E��CMH�l��YA�r}:��Z|���jB�俄+CB�y!tE�1�?߱BQ�uK
q��-YC�5�i�]�.�h�U�|����P+H�_����&�;�� ?A���J�z�
|��fv��t6�ޟ�ׄ�$?�����������|��||c�Ɵ�=�5����|h4qW�*���6�qmF	���G���/ .綍��W��	!��en��6�]y;p]�>���<]����S��ѵ�������DU� ����s02�C��g-|���p˹e�������g!l~a�p����$��;+;q�M�CqYZ������Q��ޥ�]}
��l�[VUa�5�nx��!�m�{��p������0ޟ�7\}��}£�����ۼ�/����й�7�&\}ӧQ>o!ښw!��_H���~]8���y	oY^����,�� v�|?��6�߬w�+O���T�bx�9�t�z�u���EFP��O0��
�_������`+�]����	̫Y�ζ(|�5�Gె�����꺕���� ���W���/nT���#��G|f۲B��@"y�u�W_�Ҋ:un��uX��,�ۊ&}|B��ZKs��z��#�d[��f�ڷ�!te"�5�i�XTQ�kެ�)(����Ê֍��_M�[��ҳ.BE�bu��Ek�x�
,}��Z��F1,�uK?��P���7aϞ���GԨ i��{��4+/� �c ����ވ�ͿV N	2`�X�&,Yv��P�"З,=˷6a��P��h k.܀��buݚ��������t��f1��Den4<4�|<��e�sK�MJ8"ajB}�n��&Yjʄ}�lg�	yV<C2W��	ʳ|���,[�/�t�5���J]�-}
p�Ȩ�?v��K�L��H��5!�%!b*� �[0֧���aZT�p��g�}�w�)���F2���&�	d�4&���G۴ �Z�q��'��W����hܻ;ۇ��Z(Tm�T,��Q/'�b�3w��7��Ϗ][6b[�Vc!*B:bb}JV�~���pɵ�����a�y���a�XoGGLl�Va��G�W�QQj�����҅��:4y>��H��X��=�̔pf>vo} ���q�,KK�t�#�Jl
���;�K�Gx�OD����y����i�}�ī�Y��� 
6�Vqdk�v�j<��[�%8��/z%�����)�K^��8�AA��2�%��,y`$ea$n���[/%�+q��Pd<�6�%7`��ÿ�X���d�ȽG���|$;Dw�w7(E����(��"�����&���k�Ϣעg�,<p"����ǖ��V�����}Q���`�Ǹ�^A��:�B<��]f�ym5޲���	���[î~�fbj>�_�,'�N��н��El=����w"f��OEW���y�R����M�g�Z4���[^B����Rע9Y��^=�?�_x����FF���o'W�$/��ɸ~��C��,��|�)|�YQ�w�c���w_�I�u¼)D� �b��-�1,H��#-b�/��n�}m�I�\e��
����S1-��b���w�+���؛�J~GL�[]�O]T����_��_�\�7E,�K�"GP����u���	�*���u���O����5x�X��P�Y'\��w,�Ϸ�� G�/�Y���_F�F��Tb*,}�uy�xy5n���]<���*|��P�f1Ɠ"�Đ���ը-��C�k��lӻq��A�JhWq�޾���bp������B1�I��s?|�B\/�m8�(+[�U���v1��"f1mn��o�P�va�4��u�ů 2����J) ��-E�x|uѢ����}Gā��֍G��7/ă�D���|4������GZ���m��lX��pRܱ�/�'���R������o߿D8t�O��hRN�m=��1d�C��>�����m6cT�r�b��Ou�5�h�i
��kg/~(�mȟ=2�F��P�`,%�u�~w���qyM9M���A��K���k�*/�Q�~�S�hPy��x]����hJ]IXʳ'G�	�}
!�A���^�����I��}���#quۏ�u���!E�v�u��I�>�%p3�����q�Kyݾ�(>p�a�����$�bB ��t�1-���e�Fz��!�y���`�PSf��߼�|C-���^�����Lѧ6�gO$��p��g��rC� ��>Ǯ#a��)���<���I8�"=��S�C++��.۟��Ag1�l�<|��u�'a1C�Oڦ��3mn����Z!TJI�	�Ol41����&k�i�7�"�27�sK�	�ØM��o&����/�;��9n
!I[Ǌ�!|��&�-��@���0O2C��M����芕�P��h6�q��;ѧ>����o
ꎃG�9���>�rs���4)�N� 	�\��W'ě�g�6�R�ki���k��I<�>��ӌ��ަ�(N�l��(,Y
� ���JA�S��?��]�M	��u`�у�f9V}�nV�b�(�K�c���O-��<�Z����Tr1��7���u��4�P?�s�1fF�4��V�P]~nB99j�9�"�D\�4�g�jB���p�h�|�BL_/�z?L1<�i�>�!31� �TH}ک^��Q����S>h2';'�?��L���RB�<3�^|6M!��-�G�w��<�'0�8Y]�|�DW�1Rם�&V����|�Zl�1�r�E�"�r��O�Y?��/�)��O>s�
rst�KnAϊ����969c^��]��(ׇ��a��\}�C��
!\n����H�}�twU.�&�\�^C;�<"@��F��"����tw�'sޱ�#N��g.9�f��@�f�����!������̜T݇���c"K��D�1n��y�5�$��i�N�Q;��=�S��^I�R(��Wˮ�4��J��u�=Iy�֗��M87E���644�Dr)#'cٵq�:��4�"���7d���K�:��2�! 9I�h�̈́�x�_���>+��r�ײD,������Y&S>W�O�Vݸ¿���*������9�"�%�){*���x�g@��Y��/��c��wc�]���H&x�;ߊ��K���� �^W��'k{q�]w�A��/++ŵ��>�9���5c'��p�9/R@%�n�0������s�0����AH�7.���?�H$� LĿ�������@_��=����J�Al��B���X]Bii	��[P�O O�*WK�di!P9��Dm���E\͛��d?a; ��,6�#�IB!8i�K��;��'Ї�s�g6<����E��]
��s�X*��v�8���\|��O�8h`0Ǔ[��x�I�\�
����^���$�`$U��@}�J���̿��yf��L��4���k����-7Ll|������h�r]<1RRf*�%C�`�I,��c��DLh��-�����iCi�����[<�қ1�v}����n��⊍ruOo_�o��$#z�D��'%��]V� b��!>)*�� Em� ���Y���1T�ּ1}�eSLL��1�}��]�cV�fFyY��5*V�Z��#��(��8,��!�J;P��t�ir�7�?	��.��".bӢ�5>)(�[�<7�坐C<��	A/X>��"�|�䖧2f�Ī�Y������2���C���˗�I5�e�I�,���>��#ibT�S6f�\�S��0��(�8��z��N��23m����K�8S�*�R�H�$(��d�>$������"�D��V�Àf�H����s�z�ODD�^�-P�)'l�G���R`pUy)"9�hL�)�ז5�ׇq�����P0�E�cǠ������&�p�,�nj*�8{b���ߜ�^�#� ���ڢj�n���◝�t	�Gr0��f)c~�@���}~3^���8f�����T\�zi�>�{�,+Kt�I�Q�������\�b�����񛿄����x0�=X�>�*�G�>�E!���Q��ڑ4�D))$�� ��ea|��w"�`������Ư��ʰo�L|O�?�����9C��@;�'����.�}Ǆ���b~]bb�����N&�J��ʠ[��!~���A�rJV��1���B�WU�$FOw�*�p�D��.'�ru�v~���G�1|��a�~d+�Ǭ,z�@��á*�~�|I����q�?�6���gPG�U�����)*).�֣�%3$�L�_���2�T�oSot!��B3�O�������Z�"ĺ�
9��
�D��c�L?%C���P��ʪą@��Y�ɢ�BS�_��d��sޜ���A�pL��1G��r����Ю��;�E(h�az�3�l�)�����$g ��j�V:Ru�<!2�/{c6�z��%���?��0D�O�~����$���4r�B�AX�Ō���+͘p��N�����a�ј9M�n1%�Z��a�f����b�-�5`�Y�v� ;�5a�l�oj {�?�H���9^������sވx���8v|P����Б�*��/~�Z��!;2]�P�$�I�� J������?��ؙ�"�!�8��ԩ�h��˜����b�מ2�=��Ԧ����̞d���B9/��D8��?֯_�b�!ñ6��5����� FlACc���L�k�C{�Y��p4h^��̇���'�N�,����.cbIk�U*�G�`^n���m&�A���ƺ^9�'�<[S�V��D6��>P3�{�W-���@ ��������B��v���9�^z�c�D
�ΰ�qg�o�ch�� ����	(?dCQ=���xC�B̻��S��yQ��2-��jq}�����"8��RN,'9��{tM���oR'�Q�P��a4Z%X.��^����kUb�ރb�3ڕa����#�eH�8'��9�B6Mž:�W��+zȱ:�C�DpU�[�@�����VN��m|m�h:�'�Чh���d�=��c�4��v��$�M9�h�Zu���\�Ԉ��/��M�b��S�Q��pj�5�R�Q/T�/��ADcLr� �T�6L��'SɄ_y���3��t�$�]i�PGܳoV��u7�W�s�38��rǮ�������}�oN��C�·6w��Zx���l���zm�pF���D���>q�"f=��\<l.��<�I��s�|�p��X�<��ʩ���4���F$D�)+����,�O����1�Hg� �χ=�Pk��Β	z-���M��訍_�T���:�e?�]I���x#@�S����6��g�JS���N��G���H�8Q�=a�n�������"�����m:���t˩5�(i�`��b�%!�X���Z`~�K=�ŵ���k��R�5�b�7����F {~É>}�gڔg�=#�K��&�I�H����BW���ocK��2a2%�8�0TpAA߸��ԕ+��VC� ��y����tI��n��m�c��z��n��*�H庖�Ѣ�]A�_�|��+?����=��+)�,#��ǅ�ˌ8�����cݝ_6�)l�Ϳ9����n������:���@�>)�s�8��`4�k� ����'B
w���R_�aw����2|z^����ӥ�i�p_�kꃂ�E��K�j�Εa��� ,��U����w��]��PQQ�?�)|�8�������Q����-�s����yJ���m�����&��\K$�tA�%�㐑n� >r�"�d�&50�YV]GU-�.�NUO,�,�5P�V,LS�X�GI.�B#$JC>Ya��ExA=����˔:�A?�+K����8��b5�ŕ���>~�1�.fm�p4�$��&��b�gOmc$iT��MmL=�/:�}�#2��	�'BGR��WL~�`�D�<V�|;<$@�ca�9GC1��;��:���z��dO"+>����=τ��^�F�Z����>��;�o�o�0�O��������v�����&��w�����D�ﮰ�SÝ�\����Z_$�O�߄��Ѵ����΃�zƠ�ht8z�-��;�9�vv������X\��/��	��϶��av|���l�q���;�Z��pT�S3H��Q��4Co�v�s�4��}����Ǖ��/����a�M�'�$�)=�$~(X%��hW{�a�)od ���\����ҏp��c�n:!^��Z��s*u�hg�0���-�&b���qaNu��9�\��
�{���Ԇ�i3k�ge���j<�,z
�?�RW��y�*Kh��j��A�����8�-�o*y�,�����\R��s�)d���ˢ
��֧~|C�
��3��XW$�����Y	���7���}��(
jxZ8�p�`��Ѥ�m��V���Z������+D���b��AΞK}���ۈ$m������f�����5����)�����j/
īX-�a4aco���i�Q�4��*�q��H��"b�K>��L��yȑAK))C�b��2�~�s������d ~�=tRq�{4��S�M41�n2O%��{�L��&�s�EE:�_�����E��g	#���L�	�.$qϵaC�!pk��6����zC=|(ncG��t���R��s��X���y�e�AQrHwvD�v�X�q���ɅE�mn���s����AT��{��ykX;�=�gy���s��cخ
j4T�bs���H/�O�]�(��2]Z��&��Ԍ��-:���	Ǻ"R�%D�&�!�/�)�gT ��!����&��z�==��=`_�D�ʪr�YGGt��q8	81�����7�wb}e�e�Z�h�B��	|���?��%U��/Oq��rϕI���-)4�^-DMvOJ�ab��a|�r���C��j-Q���E�g�m*����/��a�r����]A}��HSz��A���(\A��ȡ�!�A���}x�1��;��P""O��C��8�T��.�=�!���,�(s8e�tB��O0�rv��L��?���m���u7�W�De�t����~+��� ���:�Ƣy�1�i��=���z��8U�v�ݏ�<��o[�J���P���w⎧~���G�kQt�`yr�����PW�T'��Y`D�3�2A�N�Q<]\#��d��VS��Ǵb���m�	�u��y��*!��4���U�w��8r�D������h��9 s�l/|G�O��ǯ	�>�K��2�x�m�{2�E�I��w��&XPU��V�1'j^���M�5u�C�t�vFhJ���7��v�O�V=�B��WҎ	PfWH=Uʋ�pѰ��
Ȫ�E��!�4�ISe:��@�ꛓi:���8��@ �J_�	�����g3�v��椒2�<��we�݉c���ZR��[e��jqi
�@wa��h
�)��$w�j���Y�s�C@o�J��J��r�;�˰4�:s�rm�ǚ���4l��N����UY^.�k�����\g��)�U_A~��,Q\���҈��	`ѢE�$�R���=�d���k�z��\�%�O`�h��Ԝm;<��mV7��� ��v�U���ը^yeV[Jq]qI).���*,�1��9&T���q�57�yN��mC0;R����I��g��R���q��KǛF`��QYQ]�7��3J����"Y�����#l�<Vxм���Nۮ�d��w$���BZ�/]D�?I_����z�櫉�N���'��}X��G[=17�I�kb���Q�%�4c�]�m���e���H����h���6�=����f�r�U�or�{�e�!1��Cfڴc�L�[��Ox�v��NQ��SiDؙǎQsf#�S��:c:x����{�������:ӎߴ����9Ӳo�:$�!�BNe��DV:�z�C�����0�������v<�׳�� �7o��t��K3� �4�t+C�x�"��Xy#5o�|6��,�{��O�R��Jr4�.�Fj�AM-����A
�ׁ�K*cJ�znL!������m���v��F-�<{�aym<�80�N���eN�=�[���"�By��z=��ziF\�~��ě�j�/3j&�YNM�xJ�O�RW���:��L����U�kX/�G�^WU���r�d"�y�Id����c�Z;���2�
?�}p��9HL�p�'���:��Wj�^��\7��d2 �5����
a�SEH�%BXL��k�f"��D��T�DdqAhe��2+�I�Mgc�y�R΂?�yU��i��^�3D�v8	m���b�H$	�CnZ�S����'�%* ڸ���!��T,*�r�T�~�F!��)Lv9�t��\Q<�LW��ϴ���^<j�A ESxhR�\0��e����1S��~����9A��V.���uRr��iX)�&u1�Z#��)�p�ٹƴ�NE�24�u��
'͓ ��+��3�:l���C�O��y�7ݖ�D=qs&�8AV]Ѳ"Փh��/�F��I�-(d*��-m&��8��:��I����<��"���d��\q�g��,���<�$saKqs�Y�A�BΟ.�d&���{�d?&�J!k��,zL�1�\�a2�i�J#h����N�ua�m��=�Q�ٽ��r�7�Rp��A��>M���Q[���ݖ���_f*�t�S1-{�L�!i+��}V���
�i��1WO�Xw��&3I�\���1����.�ud3�uo���/�m����P4DW����XK��4ԫ��#�c�<�)N1�R�.����O��%<O�we��Rf9'"���0`)r:\�L�L2A���U7К��eG��
�暽�r᠝2qN���ɱ�������EL���x@5-[�ɯ,b����|r��7y���t�a ��}1������9f�3�s� �O���1i��Ǐ�\g�RB�E""��L.f�,Eke���=�#d2�Ho�鞛]�%_ �AJ�gˁR��"�R��ĸT�+�h�Pw<�2fyёd�Q�3���9�x~*�|
q���!S�n��CrsI���|?j��s��-,}��H#�Ф����� �>5���Q�B������wY�D�E��1j��wf�OD�bXs�*q僢6:R��E�W��4ʤ����g�L)>�V��ZG�QD��
�"A+����U[R�Mބ89����VV�q�B�v��J�SD߇���ŮO��6
�P�6;ʛ\q�<��t	q� � ǩ k��^Z����Ŗ6Ag&[{m�b�^8)���b��$b��sj)<qV)ȣb}�)��g��ٮ�B3�I��q� 㒺|����Q��:���2��L�,ۇꯡ$���c]MH]�rۨ�~0�J0S�J�����E�>�����1��j("�;b	W��s�{8+4���2EU���U���"@�}8���G�cǬu�*�E�-����e�N���>����/���<��g���PL鄩^�̳�o�dTXb��"\P��A�+��5˅�m�{ЍSqL4.X����� �PLq�Dȁ~��(�V.D�8����4�dr�\9��k6E:��I��$����3:Y:�ku�1G�QܱP�ѕѼ߯�JL�=X<d�;�1oymO$�g�Fpò"��g��$�6R�cx2z��M�)��@�&�Ϸ?@�k+D���5J�X� ,��Enp�	���B��R4E���Gt����58��XC��:Ǵ�X'���%y�8���ܱ�<U��Z��#:�}����犕��쿂1v��Ek�i�$n�D�D�p޿�&g�n���~��Jr��^���:z%A]�G�� � V(���K[H|Ur/7�<ѫ
'[��R�^0+�8p��#I�5/J"[�D^��p�]1$e�3F\����(8I�?�\�TL["��Έ�X������e�6�]�OR2p���P�:{[��}=1�U�g�`wWT=/��*"l�CQ�#q4Ct�Kh<��h�Šj	Y�ϗL���3��tp1�Ef�Cl��ܫ;䱪���ci,z���q��<YߡJ�/�m���|"Ǔb�%UM][��Ӎ#h�J�Y�)�V��:�7-�QKq�J���yb�qs�R��M���GY�ٔ��c�1Mn�G�K��s�:A�˩Nv�ɹp��i'�-�g�K1n�5�t8�w<� U��[��c8�W@J��Mм�v�SH���j�yi���\�E%9��$���Y)�O����)�2JP��y�_WN)�+.jq��Q+�a���HH<Jlڎ� ��ߦ�ټz��"f"-sm}֭,O�yΜ'F�u�rNF�Gs�Sn�#c}��ջv�N��bAE�"�"�V��wμ\<rh�Ą70�N�4u��+aE��%��<���ǡ�r�t�`�c�q�Ǘ�f��w���1|'���D�S�b�]id6��F�t"n(�#C)��y��� @����pS��G06���Ή���r�RǱ+���*�Is�C�T�O�ҁC�5|良���F�QSq�����Ն�^���S4�t4��*�	���s����Y�D���W-�w-&o���-6ƊZMkl�����|��hV�~<�C�M�M����M�N��U�&��QtȜ'Z<4�� Ԩgt��ꍕ"��^T��Z:y�-�6�q� �k�S�Җ��/�?+�v�����c�+��p��
X�9�#ӛ�$�g���Z��>v��p��L�s�T�(���o;'*H��4�nB_$���vx̤��(3��C�|M<�8���]+K�v�]by	lDFe�S�~�x弿Wt����;�MX�d�KZw|��e�'�C�&$0��<�7D𞨋 �E�(df��v�5.Ff]d9�P���1������Ds���C��&r)����V8 r6���WWW�b��Q��("��N|���V��B�3�!aE���	���(���(?�A�p�T�X����A @�p��*V�9�D9�9v����0.��shg=�΁r�� ��"�����NiN�3P<2�8��F��GM�!#r��I稩�2w���[oI "��=s��t��c���\���}'R�3�$Rw�����m�=�L�{#�#gcl��ɋ�1ǌ�K�\�&�$��r�5�?{¹9Q�CU�ND�"����8�$��㤽X���}W�s�5Ǝ����8�t��\%��;oS�P��ꓙ&��t�Cd�W�CI3�������&',+uV)��ȭܧ�;�,�$�ވ���c������6#�3M"�'|�ͪBQD�S,1Q�S&wV�Oq�Di/+�9bI��Z^�Sg� �g�jWT�F��)�B�K�T��y�������CD�sD����S!:���/�]����䲑2y��L'j0��r���L��sH��5a=���F��R�e���
*>�q!RS��/#���\�8A���f� �d.1y���u
��{Z��@�&Q
����?���1���*��v6|�)�c��9&9."���=�\��B�k]N���:?C��U_� �+�l���I��r�B���6��f��=��1��+��@�CS�������K\�Y]�E('�ͭS�[�S��Nl�8�H��!��g)T��4��A6�r^�M��8�U>g�a��T�;�˼�C4LΣ���.�r��Tnju�u^Vb��4ƨV��.�A���d�$8�x:-ST͹�N����bל$����b����F7�cE��|�Ikݼ�����&��B�l��+�^��L���$ }�T�л��^���:���"�吺ʔ���R������F�)�8c:,�צ3��I.��M"Ӧ�>':���&��?8�^���cҮ�Xu(�ܱ��@����M��Kk<��&�����2g��U���c8�\A_�B�gd7�r�/�|U�J`�j��r�CYk�:SN@��e���#��*���?a�uF�p>�r��Nv�N�2B<�Ek�J��f{��}*�J.!�Ѽe:�ܦ��2������S%�9�'�E/|Py�cps�|S@�g��	gb�WnL�e�0I��Q��4�i}����;t`��ϝF��Dz'�s*�8Y�WS,Ѭ���p�J�kEC�q3anɤ^CNbZN8�}����309����>�:��aV̳-f�f�	uE���I��.��gPQ5Itq�YGIg��M\�$��A$ЙM�M�_uu?/�6x]�+"f �5ӵ���Q�p�W���!�7��ʞDD�q�%	��8�p����� f�1%�2�43�D@.Qi�}Nu��NG9��Fky&�wv;��J�ce�i��ƴ��P~C-3�d��Y�}b'����l�>17�M�>��P-*/�}���Y��X*	U�C�a�+�G�cU���4���ݦ0��!lTv���(���'�K*���=��R>��X6���袧�T[*��Y���)3A�X��)\1d?,�a��^��,�w���0��^'���E{�#n�ZAE+�����>�vJ8�����z�7WP&S�Ӿ��R<��R_��Ϥk��<��&�TYt�Y��e���z�}�F���ey���	���5ϫ�`}��7=dL��P֩�t'2�P���0}��44ϫ��01c�1񙓝;mY'T�odx͋<�֐���)E�	^��!�v�~�e4�xf����i'nSI���!L�qvR���ʛټ��:�d�g6�}&����x/�"�N2����X��
u�N3�b�ݎ��fI�;nF��+����Dj�Y�S�c+}(W��c�Z�����,�3�����}�U���ѱ5Ь�e�����5�ډ�2KR
����I��5�:�(���LΒ��o�p0�`��NOXR�B�'�SX�o�4��Q��O��y�:�vS�B 3����ދ?�x޵�De�on�Ç�������O��޹X�>�\G���mNb�'�"�/+�W�עs$�����ZT)�?o��Ҳ�Ԏ�~��w�g�Bl�x��y�o^\��\2O!���_��>��o_Y�����ُ;^�QH���$�s�>�G�I��8�R�~�6B�^���ksp��R�r�%TV�7v�Л��w��%�[76�,�x�|�jg
�;n�܉��է�qY�Ƥ6����m�~��* ���*͔!g1�+O��޳T��
��C�L�#gy�/���ۨ�~�X.|�a�)��������}N�$s����� Mu�y'�h�y�K�:��7.��I12�0�\���o�Kp��K���o�FQVЄ[����_��ԃ821W�f�%��"4�Ǖ(��<�L��܅���Fݟ���n��m����D���W�êP���?~�"l�?��)J�)�8^O1ű'��B��_j힥����e(�ĥ�������W����w��l�,��w/���.�'M�՟��^��:���&���&6���P�߾P%��գ�0M'�����
��=�*�g"H��xa25S|X�I@���RE��3G���U9���mQ|Pg}�6����G��j]���S"2���"�&��Ay��/���:9��Ib&�Q���j22�g�7E�p̔Ɓ;�+uK���E�E��t?։{��s��~r\���M�6��x�[��M6��>�)���1��<�>Ӏn ޻o@�R��EG|�:T�����l[%Y?xpI��E?�j��������{Dq
E$�p�菜I�����JI����|*U�D�l"7�B,�o�������v��J�_�����_�E"�9A*рOOo���VP(��T�g����bi����)*�+b�Q��XS�RN?x^9^hUȾ�*{Y��cD7�N���~,���xE5��X���#��gu)>q_�B�gO����`O���l��c%	cgg����-dr�����d�"�ơ㚊�"�8R�CB���I�)��N����$���[*q��P���*��xn8n�<,CD���W��[�T	�o߿L=����̯����O=� �C��j��G���fU�N��ߥO*�|�Emh3Q9���g���˰�����7ԙ5��
���dm�/k��]W��U9�9_�����F�F�����c׿{�MM���\��nb�g^2��_D!�}��Fu�5,#�=�0g��±�:�~�_	 Y���OE]��ͬS'`���#J�(ȉ�W��LGr�i�K���i�q9	ݓ)c��o��5�
���lD֗oU�3ǭ!a�0ӎ���"ޓ<wR�x�2{�a�����٦���?<ێ��ܲ��W�s{�hVb�xm���i��3�9oOs�#uzf�T��[�55�K۸�6�w�"��$m��xjl2]sj\��M֜=SRx�V����Y4�wwG������h�09&r�L��3��YZY^9W���NS�M2Փ����~�w ��7�(<�&�Қ�\�����@��>�s�)K��[�����3ճ&S��-�p�3J��B�D�h�T�P�y�D�ԍ�v�J$�|a^1���W�+�T�����Ɯ)n�}������39#cR��BF>O���@1!-���֜����[3aA�e�)��_81��Q�b� 3z�hl>�i}p���v:B2ݓY�\�$���`��?��+sN*.a�6��^��8A���`v$�Z.�ᆚNQ,� Yv�=!��gU�T���d0&@3��Y����u���@�b���EB��Y������k6kcXf�d�;,%�X��0`N�C&�q77�2c�Il����l{�)VÊ2Mm��}9xn��F�6�-F��,�c�1�2��B��$h�{�Ddn*L�9U��L��@˄+����\��ؘ��N���f�EW��8N��`:-+"����SK��}Y���49x*y��!p	�P+�R�������csӎ���-�BB92�Y��Nuc����2�c��0�6�����lSz�[�MA�yZ(�cL�Ζ��z�Ck��&�0M�������i�\��������2��\    IEND�B`�PK   �eX�C��z �� /   images/a1fe0c5b-edee-4877-8adb-d45444225416.png|�eXU]��(��.�N�A@6�JH7�H�t�:)���n��ݍ�t7�������9׹���{�k�1�q�s-B^�(����@��T�Ah�ʆu\��q ���\ ��<����=�H�*���h��a������v�u13u2�u|c��+IAL�S���g�v��/y��_��y����PQ>~�'U�]zu��i���;�#ߐ�ʂ��!�Y�Os%�l|���1�Џ�(��7���>�So.S\N۽����o�KJ����?�H1���-9����OJ��v��^JR�e3��P��P[$�d��Պ5�F*�� <"@U��H}��:�d��E��XPF���?aF#���^6��1T�b�Z�����y���!3w��+��B|������-�S���E'$�p�մ��չ32JKO������ק���Ӭ���
���g��4t�Ɋ��c���ț���		Q�����)faem�WE��
n��������a���w�*�Ǐ�?�W��:��,/���Ζ��uH��&/��`Н�<�igZ(~�a���������ז�+��N�3w��񰱱�������������T���E}��s��s�!k4��Kɻ��<��-�0K����[j�}�5�|�,?Y��M���BLE�Ar�zqq��G^>�O���r��`�1�Du=���c��kku�Fs�������-�'~x��:��7��nnn�Z���A����!%6�	IW\O���]�}^�����Y�ҤrO15uHI	�B~F���<L_�[���xa�J��l�D}Û�����|�tbﻻ��m�AGg��������Ȏ�q�e�������޿G�DV�|�k�F��{z����=��͵�����Zh��r���Ar�ěN�]I+����}{;LSS��Z������������W����^�U��K&�	����<kk��^�1��@|&��pHk�3���O��o�$�����wc����-��Lw���+*4�ꛚ�6FsI��x)5��2����y�����DddyF�ppq�45?>����O�3���?Y"=/�{����Gܳ���c�oF���w��O���^]�mh�����>���"�̌r�g��9��f66����:cE�w
������2k��u?�
4��H��#Tpk��EͶ����V~�y�$��8�ٚR���
k��w��X��|��=
J���Bwf����2�?:���5�$}�^ԣS	OĘ�G��@�̎ w����ETT��_��質��M���T?I�Y>Ub*Wa=�(\}�� _el����$�?|�*e>��R�ڞB5�ۙ��p��^P5���_�P��E�^�/1����/��U�M�	0FA������n�����SO/�Ʒ���Ab�X߯@�=1�wJ'CLJ"��Xz�>�Gx ܡI�ſ�T��EC��k��x����6Z�)D�6!��!.(����̧H���D�b;;������mc;��)�}�|����8	7�ްs?�(��?����#'�V�B���g�8c���͚��j-x(:�fP�Ү�^:�"�D�:j����ڽ��ڃ)d��`�0K���̧��[��v��y�2D)���|ԓpE���8��D��;,���Ѱ��g�1�4���'J�1br"\`�^��@�qMe���%2�g�=������QpZ�(pY��P����Hg1�������xvp0<ङa+�Я�d�Ǡ#���v����IU������2A��t'�_���{�QZL!3���/G�
���yDP0����G�nL��b�O�`�=gޗ�H3d�Nw�X�1���$먧q ���$�NrW�F��z�+rٌ�?5j�9���g�A�X�P!�k^h�[��'��)#D��z'5y:|��J-	����h�~y9����x���(L�U$���#�ƖUW�����m*�ʧ !%���ʰ�M�W��c�������C�ٳ2�������n�T�&�R�heL|f��D��n�<�I���6Dh�����y_��Y$���V
��� ĵ0�����gX1�%[sc���y�Ijd���H�PT�9����V�&�ԧXG�{���b����8Q,��=N�Yd1"�G��EE�N��۬�n]��0���F���b����S�3M\ ��&�u}��b��ID�2�����%�}%ݜa���OX��l����QJ~��F[�Ӊ;�o��+�aF�c9�QA!����P�'C�j@�h5��S�0���D3�;��������y��7���cd��%�������p�q��׷��1,�2Oy檅��������ҧ2KF���I-AI2�+��E^!�xiiic��\M�+Z���,�� ��e�D�>/�|e�S�w)I�Y.p�i����cOϚ��4( �+8�"=���x�����eG�Y,��(R���y���EP����w��D�NBL��ht�ۅ_�����'�={FDB��œ�칒��Vm����� �۶N�������YY�Yw)�h]�����C��J�ݖ��_���>�Wt888���y��K[[��>G/��6��5�5^8uV��KN^�L^���o�.�/+��8��Y��
j�I�n!��\��\?O�/���3^~�hp :�7��>^�����s�T	�+A�4]l�~1�4Ӷ����V�Jb�EN���b��P_,�>��(		�2
-%�p�~�4�$:�)��x���#������B��-��pc��,��	2�**Ex��p߲�B�x/C
�ٯE�՝@�S�y�́o��Q6z����|EY4��A�uC1h�m�B�����������p�A�(���w
�SO��J)c�߅��*:�1�Ͷ�f;0uq�I:�2�5T���'�� (+�t�ĉ���� ��`��[���2yF�(���Ѐ�(K�E
�N�$�������DǋJq�&B[�A�z�tk༌�������`�S�s��m��%��ĸK��ъ��5�[�����;����1?��P~hs�y�I7�xQ'�%�Cݿ��*>�:M$�裝c��?��������ϡ���BM%��_��m�>X�� 
/�D�����%�Ei�=|�x ���1Q�9!#-u]p|�Ϳ�>E����f.�B-s�R��A>Ә0F�F�P�s3C��]�%�F�z�:��&���Wѵ�hjZ�%��8�W=Zi�5���Az���99y�T/��+�c�Լ���ׯ����w0Hˣa�p�����aڇ]5ޣ���s`�j�I
��m�ыLK��Q8��c��]
}G4�Z�J�*,���5������4\�B[�
��N���ڂ����k�����`��c�.�/ɐ8����E������3�F[w|O�x�`-�B�4o����&�S�w�u#N��v&l��ޣV�][��g���~�JW*��"�c>˔駄�����?�<�J
��������@fe:'�L���8��?�7pI�n��-&�3gøT端���זR"�]��}�f���X�!h�q@�1�Uv�h�~d��Pl�1���>���ī��P�b��F(��̙V��CD��Nh�q!ΐx�諯}l[��n{�{�c\
*m昦m�;E���(�'-w���$�����"N��F�$��	������\g�Ej�]�!&ѡS��Q�/D����2	�;O��m��BPM� ��/*"[�"2��^R)��tJ��7���C��A�wj�%%>�e��	|���_`�!T]?Ψt�T�*4Ę��h�:C6XY�ԧ�Vi�b�����ɠ!�g�d�V�=8��j�|	}��F�uZ�c��J)km��C�Wկ�ape��t�)��4>��>!��8��K뼡n!b�$$�s�[|lu����� �HD���F.g����R%Q	u�����'@�����1y!ϟFϿۿV�<����R"t���A\��M�yh͡8"���g��0RH��o������zdzqd���!6� ���d��-U�+�c[��~�:��=�w�MM%j_�f�H��~��g^cJ�>������Q��}���i�\�3V�9񉆬�N���:~C��a����|>�:D��~2����P���JS��ڪ;*��p���n��<������B�!k*���*YF��v�}b�=�Dj��	�#W��"`��7�-X�l���>P���&1�.p�T���AV�y��a�?Ň�gv��}�mu��/�ܾ��L�2Ě��+�b��� ��d��-U.�����ՂX�,�h��4����,PCo��m�S���mW~�%7γ���gB�Zޕ�?��1yG��zc���5*��O�w��m����\M';�Y�~
g^����	��|Nf�㙽�M[ٚ���Z=�E�H���CM�ܛÊM�s����c4Ŗ��?..����z���ʦ@���P�=�� ��	NG��,��a��_�a��٤K�0�h�*�Ϝ�j�Ԉ���U���S�a%|��H��NO�����'BY/� �����{Ľm�癟ڋ?si�60�:��~�Z�b����j���#� !��<�,d�ǽo�=~�q�eμ�?˾߉��dK����M3r�����^jX߄�hBhV�es�����l!D�K\_�r޿�E��0QL/E�c9��=89�h�F�b:���V�H�y�:u��2�f�o�7$B�=ŉ9��{lh��e��RD�v����%����/�}BC��-Nl#�,G�l9�Q�܆��!ۤ����2߲G~�7��{	T�Z0z��ʒ�x���1�x�w�D(+�_�eV� �ǝ$`�P���*����U�C>�����V����S;I�Ho~A���h�i�"V{�TA���GM;kzq_�E�8N�PF��C��6�Rez���G�C'�W[[���1��#%�GMMM&!!r-�y)���#vn�cW�$		�x>�S�1�� /[%����W��L���xrv�2���^��M]v�YGG��۟�/��$Iz�dff���j־�q�GΙ��
��'�9���
Kkz�s�8/�b�������>���տ�`T0CVsǓNr|�f���i8�>sB�n��ҳ �A���_g��)쮟�̈�oS{Kcacc��|�Cޞ��x2�gc8�����y�e?Ӄ�EFr�^���%��UuwVI��������/����"�|}3$�lhYZCHٜ�֔���<6����YxC��8LDK��D6���,�%:ZMO/[��.�����q�������(*&���˽����������s,�ZAC*8�\Vy���ǩ����5n����������DjN�ӧO������G���.��//�S1���=�p�TAU��s���X�h��Q_�@4�1�@�k��I::Uq��CD��,Ы�V�V����;�������+��{/X�%g?J���a$SH�(��t�m�J���P��HO���c�
�f�a�v���JĎ?5���*�roޔMDd$�/x����_����a���h�Ap
�e�����Q����bfO{OO��W���T<i�;�������(�&��#��fR�����Ғ=�g?F�ӌī"�DE�K�o�3�#0`�~4o�#fໝ�$B3��Z9<�(��=��Ys�dd�G���)sS�	sR�z癆���7�уD�]m߷���~2��)V�m��H$]GEv� _.S���O���D9�������W���YƢ��	0�x�'S�(ez���j��ב+�m�U��*-+���U������g��·����4��ލ���p�r���l�������Hd�G9ly(m����Q9��1�p���e���sh8mLeS���Y|*��
�Oq�x�߷��E��u^Zie�p�W��S铁E�TS*�����_�	�YG�����΅�5h���'�C�������;�%Sv�Ј�̳z6z��*:��JON�������R��vh��F������k�ږe���P�C�(��E���L���.��a����M��w��ձ.����d���h�p��(���N_D���*!!o��0�&DV�9؏�Ã�������t�9=��Q�� ��2��k����r�W0�#o�x�g� +%-'��ٙ7#jw���\�^�6��߿I�A�z�r	�z�x�|a��M�l]l�a��9��f�zk��eU��}�'����+Vݜ�[5Ե�ɕ$��		�e�M VyX����l�:��˽	@���|^��A��ΖĪuTQ���
Ł��Ρt�d�է�nD)�53���������/�B;�n�8�er8Y�̄�Ȥ�G��41
��5oVCg��Q[IY�vrkRH6mp�T�������g�d�wò������Z8�nz�M5�U�c6�Nٰ��q�]�*Z{S�H�v���Z�/��O�d:~ja���8�G�<�jd&�ci�NI��h�B7�1���>�G�򪭆���W��P�bc���3���J4�����D�
�5+���Rk�|[��KL`ٟ��dkB��:���M�y�N��%S6�>�u�<ݧ�����A> �Q�r�e
>H���7�N�n��������-�A4��Yˏ�"XP͸Zd!��3fb���u1�
0�}�c�d�H�p��u׏���xo��./��	^�M3cY�;;1=*�#{l8�������WZz,N.�cl�O���'�͓�V��[�:�^B��X�x\<[��{i�)u�\��;��y|l���a�XA�Ƿt�f1�(�_������~���Z�GVL��π-T�)w��U�*{�yz�i���//Eg���}�k�dMY�Q���*��7I���$)�X��:�"h�����2�o�n3�"�ޜz�>k�{,}Ьڴ~����	��B��n���$Ì�Jƶr������5��t�/��Ma�/�rfsC�]��ة,>�r�{s�_N�����,���I4-R᥺����ڵ2=VM�4ք#�W0w������{>�_���
�x�O#åC��y"
��;G�y����j�8�c-PTga��������/(���~_%)�j�~���d¤��vbT�������EF0yyfnn<�u]�ݏ��i899�V>�01���3KK�P�Vڌ	����$�X^K01A?~�H���U�E��ԄEHH���ǧ��i��{L�Q}��������?��4�D�A5����3�%��͙<Y��\ZZ*��<:<L����/�10��V����ҽ23#&'�`y��M�OHw�����[,\\�d��^��~�7F�~��O�ӎ��8����ۙ��)�i���@e��·�����sƏ���s˔���Imh�-�ky�eff����w~u�
H%�JQ����ٙB��)���l�. �P�4��*���@|Z��ŭ�0Z���Rv!Z����&5N�����O�����O���C$��q���[�|A>�Z^YA.{�$--0�6�;N[�<�1�/�J��xA�_eg�+��B�0߀|P=����>�*��"*JU�0��{/^�x)Yq�OKc	�n�! x�?[�ܶ������k�c{���h���� "��� lȒ���J`VV�$$$/���Fs5:�����M��i�����E� �WR2����u�Ǭ�7� �#�#�F��$�f��*�/d`�vB��X�7mC���H�-8�(~/��44R�V�z�eSᒴ(�<U����1�&i��[����'��p:(c9
sQ��}5=4�ڥyq��L������<i�S;���I�  W��D�ݸc�ˍ�
�
N..�{Ϟ?�����쌲èɷ��x�����OLyS
>c��Y����`v>�O��52�:�Y��ן_�zջ����b�CFA1<��c=��|���]�׷�c!S.�����~���\���E��ͥ�
 �_{��=x��|���D+���[W�A�����ֻ�����?}�4�
Ro�������w!�X@�a��Hz[a���F�PrWd|�OWX�����f�F}���k���P��J�Z���mRg�r��/9���x�2'�v8�PPP\�ϝ����27��F�U㴄Z�W�����3 ��`����rGXhPo��&�?�=�MG�#���S��&oo��MA�KI%k>MW����aU�1Y���]�{�am�U~EE��Ձ$�OsY{!+�����<��B����V���r�WW__��z��c��V����=@fX���$$�Z�gd|��>P(on�,.:�� �0w^�ٓ�(�nLy��	���x�}�S�$��9�<&!�Cm�ap'�~W���m�...,FR�|y���"����J�Ao[�F�بL���ֶ��5f^�H�GJ@ ���X�}���қ�߭�HQ��A�_����_n��{���	jkLb�s@Q�Oчș���C�WP�Y�������V�v���Ҩ�+���\0�(���B��Ę�F9������v;�
 �$}�B�_���1�H7cm޿�[|�,GV*'�I���=�;�� �+�+��������h�sʄ�&���־d���c�Է�X|��J�nw��(��W� �CӍ>��.$켼Yҷ�潷xp��\9砍��Oi�Hz�����)�f��~J3����*�+D��0���*��lƯUI%���r�Pq�I��C�c��$f}̙�����HFLL,m��Y���Ç1q�z�O�nt�����=zvW�e�Ս�U@x��T���s�k��^�5tn�c�����@\
vDu%���t[��lmyZ2��n�����_z��eu"��gǛ#��ҭ�/��;�oD�WV�0+˩��"�pG���8&�M�6�83cbc�&K��%|	�# d|�q�+�R����RT�|�j��ښ��lާ�*z���G%���d�u\�u$�ɑHv,�<��/<��ə�3�k٤����a��jq�mw��;��[�@<�^��*{�2��|[�J���WWՂ跋F2�/�����O�^/4 ��\w�q�$�������CR���Z��ηGz`!2�-ѽ�SP��o�x��3@V����$���S�UX��O����~�:#g$-/�{j��S�x,b� �UC%I��$AOb�bcuu�u����n��;c�E�a�m�:ď��*�F�H�� ^� �H�J
ajz6�O��2�������?�~ۥ�/��V888D��B��{Mm������"�������|��e������?�si���<�3�4ֽO�C�V���
"��;����}+FFF<��X>�ۥ�[ �ܕ�0�F��}�+�0]n9?�d4�k�#Ta�����c���s�GPAW�Õ���d�5飫��_�(��Ɍ��S|����uZ i�k�������˥C�B����yˏ$���Sj3�Yn�%�i�E��#z�,�����r�1 �no8�հ�{l��ݻw_Z��d`���*Ը�s���`5��՟����f����2���k���v��
쓭��A�7Wgf`7���f�$�ջ�	��HMe�X�G�j_`nQ����C�Da|�.�F��ԏ.�]��?��Yx9^�gі�ȏ&������h�}{�/%���"P���h��gY�t�Cʦ��M���Jm,�2%�����|)�qT�D|��vln�"�X��&��ڂÊ �ӂ2"L+-&F������_ �9�h,Ws��(�m�Ҏ۸����u��B$��������<�}�;xû��d�_bO4���9�t߁�S='^��z}q$���6�@l5����ރGf�pY�K�E^ꢖ��YY���8��kb�vZzv��Q�F�zu^a�ɗ�3:q*( $�[q�\�SG6?��g�j5�2�}�瀊���������<�������B����VD/K����"9�b*���.�{I�c����F�q)ѱ)�JE���v��ʒ���`~�,V=���l�FB%<v�T�NȤ�?��D�F
#F�qZ�eg$�pD*)1��X��� ��:;�{�Fv�+�M��6G��Ϩ���"]ѥ baaa���SE��g�؋�=�F�!��6�%�(�#�t��pɊX���(��F����G9���i�b5]�f4d�|�E�e⾾�ؓ��|�O�xԏ�%���MYed'<�FB�N�L��mEKeE���d	bbbM�
6#Y��H#�����A 7�'�[Q����Z_A����� �B��d	���J{�*U�����$[%��� [�]���M���������M�����R�����'��t��X�j�TM�� i��{���8|q�n�E%d���|{�<F]i?���ֺ�/���[����
�FЊd��А�u�\�9�<��������y�+��U���g�������81WZ=v���T��|�Z���-`@�)Q���z�����niQ�
���T�/�]*��X��#O�Β�w�17E��&*�@i�yN���1���M��� �R/O�4 �ټ9[�oԁ��Β�T<=k����\�zoo��'�{.cO7x=���k,��M�1�u�Y�n��W U�DFJ*���Ӈ�T���qS^ �a�,���
.�f�:pԮ%�nM�C����S}��$�hl9��V��Ѐ��3vs:ٞ�x�����5K��ʊ\��=I�I�M�Ա��d�b!���B�n��n��:������?Nڗ�F#��"��=i�u�ptt4y�����8'��ۓ1�U��ocVf},z��eU���+e�	7�P�<`���{}Ga0`E^�Mp�	�����o�w*�3���cB�UF�Ÿ;8�v���ly����9�@r��Q
��(;�M��oLb�x�`Ttb"�-�S䫤Suˀ#���!�,���t�k:OHjD�9\v���1ȫ�Rhh(lK%��)���yM9 ��8AR�s��~�;�_�f��v����C�k��x�I�Al��}	P"7�4S�?�ӷh[X0�����.(z�KUM젲l&v=�7�'�x��P7���Υ�U�����L�|�x����?.���s+�Ȼ���Ks���Ms��a%�|����`&7#�����`%TcО�|k�8> W+?�`e�B(g�����Y�r\LLWk��۫���n������j��cS*k��� �QVg�9����2!ȅa��aK���ܗ���2�"3��������Tw
Y�v{{{��,uˠ�U�͙�,���ny�J��t@��Z/�`v�1�V��]��,M/����Tl�;H"� ua�@]��l����V� �-����U?9�����H���^`�a���"�$�~�����U��r��;^��<z��o2�1��p׉Yːr�C6(�=F�A��5��(TW!b>���#A�Ъ�0]_)`e�����x�k.j_A���-�~�֗&z�<�ٞo���#��^,wX���,�R������~a�F���{�ۖ��_6�$+��2)@lMSeY�r@��)�]�>�u �*+k�gg'����k�N�l���VS�YX�<����F�3d1Ns��ACCC���BV���}����D���1*���h�i�P�;�r��z������o;ee�x���7E>�Լ�sA���b载���M���(���]�W ���e*\�XXP?Iw5�exuuu �\�uu���j@�����4Y̌7.�1h�IKcA���Ix��O}���BZ$���5������OҼӫ?����e~,a@V�9QV��.�WW�o�ަ�pi�\̣a��4���I&.4����'�}�� 2�����l��3Œ�3�:yvd��2~��x;�P2::��ֆ7��S|���T����k�օ����V���#ȃ��ә4��9����>.n�ˀ��e7(-����d�R��g>�_�X�Dx@�(���˽���B��J)�S�g�4@�i�Є��܊����=�茻R�_z�x�j?SE����:K\��!ZI�@��%>��py�I�_Fg��2�p~�M��
��b���KeV���X���t���i?�-Wa��n\
n�sP�a��T�B��P몪�\��E(+)����Ңc�⫠˚�kKK4�����j�Ik|5H��u�4����Yb�G3T��Dn���рY��n�+�d0�-��6u��$`�-�fȟs�4{��q�����V����gۢoK����
}����7Vvv���������{�̞{^�ut�}o�G�Җ�I8�����A�z���o@�P��p�PSS�z�n$�{}��LdA�ƆӢ���yo��'ȭA>[���o#Ș����f'U��"�5^8��ʈ|�%�3%�mw��*T���kh8��R�eJ~���%�ׯ"���&�z{�$OF5 <��ބ�R>USW��.k�?�s~�����t��O����\��&��C"b�wb.k�`�[?����G��SJ'���I]��K���s+$�/����d}`I� �n��XOO�s�&D�$@z_��s0�˗�.�OLĀ���86GH���<�3VV��m
�";//E2b�܆�����t�ߥE�hkS�6]9@�]C�
f=q<e�Fu��b�Վ��I�N�<H���=����=�J9���T���Q�롵��o#gg���.�3c����y�s�r�]�����/6br�{�;%A�!���� �TGH[қ;H��c�*'/�2+�'C���Sp	qՓ�����YA��*����%T)�@i�ȵ�c��q��I�ˁD��BSHTq�f�yO4p4�*���"�$�X�~�o�+�kpW�J�*٤ZM+���w���ՙYn�kg"����=£��k<&٭]g0S�Y�p�x���!jn���p�����t�q��@d���vb�k�ɬc���[P,i,������qD�Fb����[�k	))z�b���z�j�x<�#��w??`��}���)|վvu)-�W�ӕ����	��Fx��YY��S�z/K�zj��\��JD�ԗ�����ි�J2�0\XQ�����.x5Yb�1Q���'С@�ִ=���%��e�;4�P��쭣���J�E|�*]8ٚ�R���e���W�F6�;
ڝ��N����[��d@������a���U�m��3J{��LQLP�H��B�>ۍ��w2�V}t����o#�����q �r�#��-��<|q223C�	����齆�$�����g>�9ֈ�f�����[l=��*с��U_�$�(2_�DfBږN����{
	�t���/$�.v����9�~P� ��z-Õ-�k�C_�㣕��Tυ�	�C�%	�?I���m�}~��=1c�7oU�?���R��o�7j��_�<�w	���`��E���ϣ�c�`A����h-�؄�WLN�NmĔ=MAs��%T��4�Iȁ�-5�$ʾ�����H���Cd� ��*'�]j�qr�$3g,{�R�5���X�O�5����|����|	se��!l��oc���򗧻s��䔾a���~zt�e����`�'�/dN���)"�����뛈c�Ǐ�F�㞏������LYg���.hz0[벾����ܼl?!!᫘�}�s���fQQ*@H��>��cU��u��.�����3R�p�ud�?�I�2�;�O��p_`��_߆�}d���8\7!���� �v�W�[.��|�&����Ԇ����K��_K&!��ďD5���G[�A��"O~��"&%e����t�D����%%5��p��0�C�cPPX馫x�
t$xma����)�:M�&6j��={�IsSN3!ȋj�bY��R��>��[q�� ���r�Wqy���qV�1������y�0z<)��1+xdf���Wj��H�N����x)^�0�,��U@L2@ ��	үW�E��lB4�UBh�l_��/�g��H�����C6��� ���,�����9F�J�{�Wk}�SF�-��U�o~+�#���C �|9]a��..���rl:���g\ZZ��qf5�;�Z�ݙ�N�؛.L�����&�o�cӻ�b>�׶>cO��fk~P!٪��	9(��v/@�
��]]|I��b_�S��>�?6����=��D�G�O!{���h��ځH���3�y{��s�>:OM˩ư���|��-�p� J�p^F�>ݶv�j���ﮨs���B �Mw�,��tgF����߫��㒿WW�	tṔ`�"kc�w�mh��Q�$,dbb��jB�[��@�]��ZT�T�1S�üW����B>���4��=&x�8o�|<㼂�Vx���x���u�f�SEEŒoA,�����/:�R7�n�[����>Oe�J")�� �P���l��k��9H �Da�d��!��~��?�NK	��"�ľs}w��Gޟ�6:P�Iy0|��f�ۮ*[n���#///<���E�v'�Qz>KA��u�"�4`vXXX-�s�?���X���o�����<��h-4h�P�9��N+*)�ֱ��C/%��x�zW˓��ޅ��BtpSD���n�OC��
�>�H�9�u�%.����U�����缼�pc���rs��XI}�S�xDqQ�������s�av�'��_�%~�ʎS�ِ[.�.&�'������hv���r=��٩an^n��ACZ`���P8��r�VO����[�����|�p_�L\J^݆j)�Y垊ѣk��������Xܪ̔L|��RU��̀�kij�pp(�����ڷ��/���?K���Z�;��å$#��c����<d�Ovߙ�2.AH����NUy:Sng��>I��pZY�T��#��v�>�Q!�\��1		8f�����v�c3��H�o@.�����F��]���.4�vHި�1�E�pW���l]�  y,������I&����&�)?� S���Wn�ᝋ^������g�4�C ���S����y���	�}~hOQ���������������B���{�6m럹@0�l�����k�d�ӐQR�zo��p� (�X���E�����6**���B>�#��_�ձ�/���W���g�L���u�Sj2���V��<�8D�<��uԨ��J����
�#OA.�l�t9�T�)��f�{�~�F�GnO�'˷;�Q�3OxZ�Eoq��h��g@p�S���Eu
8}`�=�P�^����C�
�# t������Hz��


aYe���R?��1K�n|��	�k�V�|��h�P<3�
pn�*�љ����	33�n�U���;����}�w�[��"Z���wr����	Z:�(%�x�MWه�
��S� �m_�YXX�Mvf��l�s�J*��XX0�Ҕ/la&\��@�=:��|���@�>+K�ۖv���D�t�w����3��:��j*U�ۨN��! �@�f���>tߝi�@B������ BF��ˆ�~�(��9ggg��W�F��'��_��!����bx���}ΪjZ��hi�.��(v�x������3��Me�OMM�%h�&���鯱���dUX=�����L�����שee�*�ҁ�����	�e
j���	�w����t`j[Q��ii�(iL����v��a.Pҿ��.#p���w����L��ȉoV�05uP1w�)����?ܶ��^�״�pK�ӊ�����s�����/\��7Y�߱�V�ud��V�as$���W����F���!h��2�fvlfv�f�Kx��Tf�aT�;/���lӱ>�����3~���4O
3n�/(��9J9
��7�gB[��
%��Q�q���P�;��x�Ļ���x,-/h%eF_��J߬>k8��I���?)P���ЩgVV9a!!�g�s���V�ޓ�׶�l+H(2�����,�m�Eߛn�*����0Y��:��!Ec�&&kS��".m��@3��'`����������.'o�zd������!�չ�h���]i-�88���66�f=���]s��W2�F'��X��
�H��q�F@�q�[���W���%D?�..�D(�m�_�qn�%H ������6�&a����VϬ���JA��Gto��k
�;aC�O�Ɔ�Z��h��]0�4�<�'�F�ܯϝf����l EJ�j�)A��*�WŠO6x�[)�¾?������@}jj������'3 x�=|�{�j5w��_�`s��m3���� ���y̨XZs��a�K��t�d{MO�i�ݚ!X��Ef��c//1a�I���Í>S�����su�HHI� ��<��9����)*B���O�d�;&vߞd���2C>&�)���{vW<-=��y�I�(�64�%���˯EӀ5B�А���X���O~ڡ��^��&d� Nu��#�8��VV̒ny^hk�'A86�0�`��`%�YT��ښsܿ9�ё�
"y�r��`R��QP�T���?H��k���鏹d�r�m�`{��>;�U[��s��9��y:���}G���:m��az7C!��;?�,;��f{R ї�3P�
�~�u��N
ŷ���	#phO�tR�K�1�Y�D��#����tN�����+!f{%��.L'�@k����Lz�ڠ-���~1���=$��$%/;�W��y@�T���B��>g�o~c���M�w��d�qf�X?�!�,�=��?x�&K�]�ܘW!��:�Y��x;����b����Xv�%mxX]�s��Ǡ*|�7A�V�������(235f���� ׋����%]��	Y�ga��.*��4y�����&���n��w�4�����j4����~ ��Ӈ�JKK���9v���<8�X}^xGBV��iNUܪ�U�����������}�j(-��6Z�G��R+�%�{r��F��Z�;c:&n�XY.�����ic���*D��������VV�Ib~W�z^��~E)�ǂ��������4M�[퉷����Pz0M>l�(AZ�*;�d��~�{Y���&�_n�!_����e���[��D�c�fll��v,=��d	X�`����o�<���t[*�1d���Y{��R� }���%�ďUY]�踸'��ȷ��o�AZ\
n������� �ji�=RR������n�.�C�S@D��DD��Ni��.�����~���Aϳq��̼��ϼ3{�6����J��E��m�,Q�绯fN=@G�hjj�(�����p�'-1nɀ����f������(~B̍��U��;�Z\�̙:�]��mi��,;Z�Gc�Q�7(�g^Q
�ys�gy�]#ystSV0���7�C�9I�����·*�%slv*��g>��Dت������6�!�;NUO/2�E�y�яru�vp��T>3\sl�����4��r�a4+�LQ�B-yeeL��CɁT�a&����$^;bh.�+��Ԩ�RE���i��HH���/	�p�Wcĺ���=L�ؑ -�Ï;LT��O\<��E~y##��
�TmflRR�XS0LS%���ښ�@�2I�R��\ӵ�JO�V˕)jV���,��gX͍�7I�ɩr8if�ύ�/���gfw�fppqq-0;###���.t����?��'H����/��#Y�Qb?߰9SYh�U�Z걕�H����qk��v�����nv �z��������4*�^*(t�dK�[�W����>�Js^{�Ā���E����ԯh�C ��g�A�|�qh2��Z]��*��^����L�E}��q1S ^+N hu�TZ��4���S���3�'/�<����C�YdM�ڠ���a��ݭ�:���GMJY.���6V9��i��e�m��FdT��F�����w՛)ʅ�]���\^�]�n �@UQ����R�	`�W��ݑ ����cbD��jjR�##�f\�����TU���v�A����RΜ������U��>����\����t	��s�Y���k�s 4t+,P�N7A&{5��Cm;���n����H���-ׯ_���۳M�����W���i�l�Xu/3K��s%�NA+
�_���<�W����Z�]���ϯ�����U��<��Bk;�\��a�	�EY��[n:�����~�K5��rL�="c����7P��Ƿo055yy�X`��G@�wnO^?-�0�H/7�C��B��6m��J'���Նn�k���Ȗk��P7�W���G�����7�'&z���ǡ��rXl�,o@G��O��yO��CK����k:0p��[�w���

��}u[�~����} �����oL\JNI���u?T9ԋx�Jlll��A������6�v�Q4�R^`��JK#�
���:����;�{_�w(�(�����^��Epuu��ꉡ�q�}���c�c&LX���P	;�)@K� ���9���,l��Gd��B[P��a��u�ٿ��JHH@S�#%�|3Y��@�_���S7W�՗��cg�R��;99j�A���E����)�V��)�J�Zs��/۠�"��T!�S���v5^��	�Dv[�kB�����g����I!��ܹ�$�$� T�'8�X;��t�|���s����c�]�?�����s�8Z����'��=ʇr���'<��S�'qe��ۆ��^��0�����L���rb!�F?�Ǟ��h��A�=R!���6������?~�QTĀG@ i<8����,���&~NN6>>b�r8�����y-F?�P��d_�z]�����=`h)Yَ�E
�tLB6�F秠w�GF��ϖ76���9J��2B���m��$���oJy5AoAd���&���ЏD�q�V'��?�G�"X�N���Ԙt��}������g�:�V$��=��8 ��/��|��?���'K���}��}�+`� �].yl&�8x����#dM�M�Ͻ��eL�>>�^�%�v<� Ԕ��򦶇�������5+99����^��v����%E�֣�o:�"�:u42pҽ=��K+<2	�F����&wP�1����N�?G���o�����o:�`Np� �����C�����щ/���c/��'+���~��ĩ�R�al���U�r��=����~���'\�ǡ�Y���/q��v;?�y��Ӿ�o;>��g1��[(%,%���N���٩�H������|���N!zuۙ4��DI���~>=b�3e�Q��Z����'ay����V�E���N�܇$+:�[�R���;K������P��ow����f������E����Oel�Ҩ�q���x�=�X�#���?|g9��eF��}�����q�^��mh.��3�U��K�?��v{]��dD�m�/�.N{�F���� ��n��T����>�o��>g���5U������C�L��/��s8��f�Dc�Vr��3�����1[A֜��n�#Ƀ���>�s{�_i�o�yld��WE_�=���G��YŪ%�h�o~VK�a{���'!�p��sX�an$�M��q�|>��}�`v�z���HC����#t����Uэ�{�_D�k�Lgu����n�q��z���?<u�+�8�~J��� ��M�W}�x��T�Y̖-�W�$�C��级's�zt5AEO����f��4!^6b:6�\�HS�(��Uv5Fz>mQc~��}�+j�y����C:%����_;�EL/�l(Nt_�X3���[2��(Di�	�%���	���nj�c��Q�kͻ~�y�1��� {����4�'���g�ft�8�&V~XiZg&Gъgq��Ͱ�SN���N"���{��X�m�ׯ7�3�)"6�D�����9&o�ꅺ�!��2�<�΍�@$|�>ͅ������4��~��'o,�E&BZ�'Ǳ��2J�i6���#��>ޢ��b|���ll�{��)�.��>��h6%������Ǌ.�9�.hx3�x<{�^J'or}�j�R��Vr4�}���c�Y	n�#ƭ�36��G�LGD��@��U���2~��ab��j�<���gI�k�ҍpp��}ɹfO���+��D���;ׁ�jb$���.}?�xqխ/B|q8q�q]�u? �곂����[�G-I�x"�OlΞd����R�8 �CA�
�{
d�t�;�ES����1 ���/g��#�|&��̰aǅ�c���f��2�����]�Z}�ݮ�c�AP,PEL{;�h>��[fΩ�l��e�Z����m�I��3��J��� ��->� ~��<uα��S����r�z�7����|b�U��>�����8�]��)��]��[&V{���Cn���tnW����3j$�!b�Dy�ށ��y����^J��p�N_�'9�W_F�AW���t9�ɊҢ�/�i#�Cy���A���ݔa���x�vq�����b���_�G�����vh�A�f��'\�}�[="T]�h��78�Ȝ��H㺛�F�)B�"|��>��y,�M��}py���1��4�����I�[Ej� 8�`r{���s������o��o�/̳m^\ʲ̚l���L�vWd�v��<��1,���kx���\��o��O�뮅*�R�[F��c����ulݩՋP�JҢ�(�ώR�=��wML%,�푁_�.�SHj�M-�!�w��M�q[X:s�Fi-�E]�P����32n)�z�X��Yy��P�:������ђ{L�$��DSF"1�~pK$�݊#���u>ҏrr?o���b�v�*�_�!zd�Ԍ��lU���>'�]%���`}������p�5!DX��������_����"�~�� v��d�md�F�U_�L������'�F`��_��H03�YԻÁWb����R�N����a�$��w�/�&�y�7Q"�.TT��T�	�mjac�>��[ͷ,U�?�s�iy�����@#�)MA���y_B>��w���ѝ&�+������k{��[x�G$��!���uvKy��l|�H�����QÈ'vy�Sz���X�i�s��ck�&;V�iH��^h�˫E�x�÷����J�%��bonP]����/���H��]�ݓ<�}��L��8�_���&�	��!���Y*���x3)�O}u70i9��[�`B��Ox]3��S+1���,,�W���K���'f�'z�N��;�����o�ʜ80jzt�0vط�U����!!��X���^����ş����>�~��,�����w��"B����m���?���2���u��u��4;x���h��+݌�YOc%�;��OSI�x�?}�6�G�2�L/�O�s�>��uu���]�a��n�}pt����P>��K?l�Ai�f�u�bL��2XLۇ�9�9�a��>��c�y��-wʤBN�o�1�0u�c�'�&?���1_H��;�xC"��8ߏ�7h8�'���o���a6o-���Y� �=n���Xk��B��qz��V{ݫ�������;��t�e�T���*B�����?xT��D"����s�s���Xv ��iF�CW-`ֿCҿVnI5H4��յՂ��c"5Y�=�r��|�x�Je��T)�t�T1&�k#vw:���:�s���f�zs{w�/V4u��r���s��Z�a4G��
���S�9\_L�����b�?����C�wg*q�����7�?��ľX�6m��k��S �Dn�(�	��g���J��qI8}�q#�)R��t['�5�Q��m���
"�\�6�r��~�NF��
�-��AL��{꥙� �K�wѧ4q8����"�iC$Ǚ%juY�>)))#����}����qr���@r|�����!���4���r��b��g�3Hag����	�*��ғ�bC�;g^I���GS[�jjjm�{�:�O�+g>�<�H��'��~'C�䭭}��w<W
UHHK����.H:���44Sǡlmm]&E~:�����M�4!wL!�ddg�������$Á� ��~jèU'� �:�G`���	2��O�>9M	�*����2��ax��~��x����M�8kܓP(y����p1m�7"FM��G���.3�����-���ߢ���,Mf�fG4f�rߛĴ�����)���͆�/x>F@@�����\����.,|<[� ����������
%K�(K���<0������ޟj`VωIH���:��7�ӭw��Ѹ/�:G�*���rs��%�ɰ���z�!L�qm}}�z�޸��K˙�D�������KJ�à�sB
�=vQ��J��р�E�3/��Y٣ᘏ���3����r�-�O����Ώ�kϗ��P�(�Lj��υ.F�b����yk���A�k�뙚U���S����b�����[Q�!ZA���G������R�@��3�_�� �1�9�ʓu��Ņ��&�uV�-3�D.��v�́t��(��ֵ?���g��_�4¼H#����w�:Ӎ����rrs���B%t\�Evvv����떑���RH�s�hy�=Nl�����2B���UW�p\䑢�ڵ�����}N���a�^R

	eO��W�]w6������=�p�|/��^�lC�(��B{��U�R������K )*���.kM��l?���XS���A��--d��$T��<V���F�-��bk�=hK|#|>mn�,��v�'�/D��qoo��lR?{j�ܴ*�trrJ;���nց�RhZcO��%l�l��Ĥ�vvx��ȕ ݐ6m}}=��'��-�����'�B"[���O�|d�����3�oǖ����߿�G�|���u;���KIK/���w���͹/��b�e����K�V@�k��8�p����l�7&,8�H�$c
㺂Ȓ n�����|o��]������ajvv��s�/l����|�)<���L��Z6�Mj�h�3R홱%+���G���q�%ڏ�R��<A���~�:\���Z��۷��P��2��VFa�z;Y	пk��>^�:��Y����W�!I^��������GR��'cq4��]OuLLL���<O�@�kM�0��a�aa�|�g�5��ϒ#��h/���D����)S?==��i��~>��ګ����=]�ǝȂ�r8CZG'q�*Vq����G}���A�6z��Ϗ�[`�+Ɉ��7}��������Gs8Y��JI��!Ï�����X�IV�Q��ܴF���لN�YZ�$�-�ʅ]���e����C��I�x��.��UzV"�'�Dn!L��YnO@�����ev&%�8����rR~�����V��ZmE�BT��w��kt��cS\�)����, w������L���G��ۯ��M������>�R�I�����q�>UUq��<�۝.G��c��TB	����B�k��������8[�\}_�rI�2v��뫨`�{��=�pq�}�?xh7+w�����4ɟ�o����������&f`:@^����+|dk:���x�p��wf�8�V$2Z\T��:�����٨�ze��PS����ٴ�������%�tpٿB����۬��
	�^�6�l����3`M�Y����*vq`��˫���g4^�M����1
=�p��I���������cf�@#�g�6�<�O� �O �G���P�p����@B���9�\�e�5��Ԕ8ʵ���.lD[�7�;�N�5w��}Gy H��J�p�@�]@l���(뱶�>MV�!pF����V��?���(	n��)�c2�����͒���o��{|&Y����/�bQ\������	�Qg�h�d� � B���F�ELǾ����y�JE+�N���&Q�WBu������ם����?@(�p'� |�C�oOF�L���j|�av� ��=�#�o(P��4#}oΏȐ��\�t�h����$ )heǞ�!-R�R��HK�'�&�F3�����pO�������~��G�
�PP��'�p����5�z|RD�y�B�2��0��f����H1���������BB���	�q�$��/w��O��O����Q�D�-(�@U2�kkhh��,,�%u�@��'�d��i�2h�|>. +[�5!|,�($Ю���pXЦ�!��!t7�����t������ j:�T�v���%��>I4�Sjd,Ԗͩr}�h�h�35��$��'o3zޖ�T�����&�<)�j�L
ȋ>�΄3yɭ�#-�΍��<��(��$B�����i6Ixm��x��F��D�+�hGA��dX,�c9@�sQ���}i�=.3������*#��>�mؾ�g�O�=$�HȂ2��.�Ӌ���V86B��`�C���}��s<W@� :�V�N�Zm߃�$71���� j�D�8ߝM����WWWcGuI<'�p�f��ύt���/��-�� >��L]hT�2�-/	�^"^���n��Dϩ:u�ҳ�Ca?t�p9=?�O�X	7'�#�����CCMM����Q�vp@�������U� ����geg?z�䉣�5��J�a�@�x 9��LP<>�4� Zr<�Ģ���3�R��1Hq�����q4DDDKy�a�T���ttti�}������			���k�0���&o�ݯ:\T�H}kC�g���ĸ�@�Odh���4���qz�+gF���]���G��:/��2�蕼�y��B�	V�0(˅4���Ẋ��������`df^ٽ�}������jh�e9����*���?�|>*''���yBKg9�!c���(��h�;�c�~�����i[ޯo�E��"##�0�n_.����R�u �q�E8�z���Ȯ�t8������Y�)�����8&I�%<
rӑ��� �Z�}Q��	�ם���_P�b�|�kcVWW� 1����vO�NL �`�oi��;כ��.;�C�
�92���o����,���l}[��+��
��Z�9��N�8�����w8�,p�����{@��W��R)��9���0�Y��CB���G��@�S��,��;½�|fVNę�0�{� �i|+d�����yFF�V,�KɁ���0h6���L��g�?���>v���|$���.���KG��WE����X��Jȧ��		e!�S �%G{�Tp�ȿ��oR9�Uϝ���C^�b��QPdfC���!�:�t��ccc�n��ݙJH]��l(��ՉS��#�Cawޞ?]�A�-q�]t����b�o����.vgK��
O@�[]�t�����IB��)�71�2��Q�lUJjj��Q-�t��(�Y��E]߽ˮ�M�-��&#�q~�O�.+H�0`ٜ��2�P�n`^-7��$;U��ij�b�kA���Uk���X��6�p�h��ugF|�Ξ&&T0R�6B��ǂ���F�/@���߷���b�x�^YY���1]�o�h�`�d�6��(����c���NЁ#�����_��d8��B������S�]�ؔA���Yx�����		]�P��<� �q��L�;���J]�%4���ݠ��+�QP`5�D��D����? 
�������e}�WB�����g�^�ܠ��̞���iU�n�Gm�)� �(�ˤ9���'//��MF��.+�$Ez0�5V�@��灈�
�GIIMU��zC%�+̜��a1gS'�+���i(��?4!�q�� d!�CJ///~�R�����~�����������S��;��������H�l���{tt�ʜ 7������7n'	�舸�$@zi"�_&�N��㣯t����}�\�a<�*#�j�� X6хW���V*U�4� Ã��CNxYXX<_����AaceuHD�M݆b��\O
�����c/[+4/��ϲr���3�� ��|��Ir�j�&HG)0v��s[h�aNNP���s�ǫi�і#��4ff4�M888xxi� :s�Y$JnS$���ÓV��Յ��gi`@
�����	����l����r"d@*�=���@9� Q������H���W\[��l9�~����@>w�G��_456�S���0�ɡ�>���ɁA���٘>���r�&z3���E��`l�C�o��tMV�߇{����O����lQT��"m�vb��k�M��Z1���(��`c^��O�)I��x{{h��L���b^��8�!���򧤤�F�"&���S\__�cEH%%m�
�|l��������s���BE6����Q�޷��� GĊl��5@������9��Ȧ���TⰢ�;cK̍V�oʙ?��K��e�6 ��5�j= eb��kg� E���&��2~*DDH�		�|0t"�А��5џ�M_@��F6�z�����		+i�1:L�<��|--ݠe[�Y����݊����������?ha�Y�V� G���U@9"d@m����D��C�߶�\O�xސ,ǈO�]()�-��G�2�lE[V�gw�T!��/Y��z�{���G��CMO�f��F>�g�� 7H��贮+�Ȅ�8�s9.I([r`D缭փ��s�؏� m���ưe�c8�j ������NO뺡󂬗;���	��́z�['X*""��g�V�7 �ĥ���lT.�?�4{ LPPf���\�CҴnJ!m\\�n�6���ϛ}�[��n��!�15�6k�e�"M�_.~�, ě���+3ib�gL��N�aPN���7#Q23�*2���v'-ɭW����R��ʦ�&�v5��@�q �߂DfZ�7:9�����^���_�ek�f��5C��ԂD%���?Pn�5���I�e����#�b��qR��*��}�ǂ	�8�&�k���LCO�:[�ًJ\�ޡ��������U?�@ A'd�[�;�z[�n�۱�
B^�E��%
��$������ߋ����F���h�&����mu�7�WA���ϟ?S��z���b�V���cu�Y4 6����>m�a(-�ub�E��x\�'&&t+�<!����7�J�[wHቒQ�L ?�W���׵<Ϩ��`�R�$'�z:����B,�ᘵ�':::�Ga�|�������Ǟ��v���ms�5�����~̴�*��5�C�0�􆇃�Ӏܣ����d��S�]�)DIsϕ�^ԉDh�T�r��(==}�����Z��d�8%Q-}�vq�X�B���}��^@l�xğ K@�����BLi}��Cy�֫&��Wkx�b]ƌ1������@���R��w��d���W�64���焄�y:n�'41�}��r@5`��0���eCV�:g5g����ޟXɅ�Tgh8������G82*J6���ƦX�o�@��0_�tk,�q+�.�^Fc"%E愕_,��_���[\�fr,�ꕜE�z���7'����!�E���	q�7���t�48??����d��\�6�Y�	�����UUU�n4�
���񥅕� L���N%$|\�-����T�k[��7ȞQ�����ς��6!p�p_%�in&�$;.N�����MR�i�U�&n��"��N��]��|d�:9��!Z�k������ݻw�"��i��B����w�-� S�?Q���k��k�`E�]Gs�����F��dI@�bb���<���nv��%����n �������v��'��f���?��[�d��+g���:e���E��޾��Y��pp(�)�.>�������e`�Ԙ773���O|����m��W���B�:#>�z%2RR���O�=�l�E$���o����G�Ѥ��:�͎���0�o�Ɵ*I{�:�m�+�_�psts �V�+<k{�c����lk�g���C�L���^�ax���o�		�N\E��߿c0'DF�D�5___�,�� �r��_I;�^�H�����YUU�E�Qb>˯�wY��&����$���f���8�3��K_׾8W�w�v1TpG*��!?.������~>�_�s�Ż?\|���>H_P��{)�9���,,�~����wa�С.�<r��<l	��@� (0 ���1驱����=�hF�|u�]{nb�ɹe�V+�
��Y����6+n���[�pL�y�Jf{k��qXu�N���q�\|�V�<�˗/9�0 ���݄`;��_�� ���r�o���b��K��������b~�vvv ؄�S�[X���� Ϙ�+����o&0�(�Wf� -~��-��Hbr���4�ػ���x��*��d�#o;�a �Bs\ #�j�uk�, �����& �|RrUИ�FzN��0(��, ̍x��T�YQ]f�b��QS��F(��Ҕ7��g-8����0Ã��@3�6fm$9%(r��մ��݉X���֪xF:��`5�+��N��:
����_' ��WPP��{qg�ޅ���B�?��'F�L��Ё����j��X $�P�Ѯ�B�Й�*þ���������頳WKm�܄����O��f��T�#�I���n@�R32�װb
s�^G�����薫3y���i�"�J'�H���O��_�V^OTt�8��b�����o�@Tg�T@⚳@���*�xxe��]��E����%��O��cc��!�N!A� �CU%�?ϴ�%�CǷ�����=1�KMJ0�C�?U�Ry�Y��+�f�%���֏�� H���A�^�ϭ�L&@��̰���m���d�� 9P���C�l��[���ٝ%�S<}*�zM�l̷��ͭ�#k|�����u��_���666��+��fs<W���/��c
�˛��>������d�%��g6�~�~^S��(����@i)�:��vp`'&&��&$#�o̬���z��Q;d2��o+n�o��=��>���I��}�2�g�**ßk��#�������ʏ����ӧ���]��؈P�-]r�`�L�O �P�ũ;�_��2��������}H��N�%����(S ��{���~
���A��ҲhN�ҌA�L�|���8���hy��S0Y�Z��`o_�[dH,��q�YW��uE�����&����>/n%]����jf�&���x}������:.�f��oѿ����R�ZG}�3K�ү�4�'������ܩ�0� ���z_8��+���U��x���˴y���`o�u�O�b�&Z�Ķ·�W0ld*�q�zT����x�k�b�{P����j����8�j�!P|��q�=TXf���rA��*��p�i����g4�Z9gK����&Wi��`���&4�H�g�F�/�k@�m�	~B%�4bb=1�?��B~�i��m�]5|����\}�* �ibz,Z*b����E����뇱����憆��M�bI�Q���C.%7	�^"�q�����ђ|�g�]�P+�oS���������IO���L��3�����)�JF���U����#/G�xI���\L-���䎮�i7O�jFH�0�#8��PᆞO���Ѧ�;�R����_Fk�rW�=����E ��D��h0�t���ý������7�E��<�_��:	��t-F�>7C�m�Z��jA�;���R�L�cT�����w64ד �6ѭPԘT���988c*^^m�B(�ʓ�#M��"s�Q�:�ڃ�m+�n��ł��k���ݔ��A�y���e&!%�S?0��WX�R_�il�TK��Z�+��[K���}Hpٕ�|�]�ϯ�]����"כ�u�;�bl�N�oZŇ �ߐ�|%2���1t�]NMO�GB'��*12�2���s��o��l��A��ښ� Ӑ������������rK����Q��Q �1�aaaL�D}��S�憶q?&!����=AF �=m-�D��F	���ԗ���{g3��%��%����LF�n���.���Hww*62���nO20"~ �On|j߸���L�w=����aS�"/�r�bhH����q���x�� �w�IGy�ߣg��C�T��
��l�X��H�:�ez[I�x'�aG�I�j�L�Ӹ�𨩥�^��$ccc�ü�J�<�[t�Q��po1_f�`_�Nට���r��t�M",K@$��⫻���3j��><�z�x��d�����S����ם�i��KRT��'���[Zm�ya�0/������u��;y����i����
����~W�89���&80�drddda�B=*�5��l���_��a���s���˦���W
X�q�PV.�V��͸q#B�Q�k�� ����KjiM$��4�9����1t����INJz_m3v�8�D����7��\ۅ[��Y�GI �}������W���I1m�����q/fǚ�0���2-�ttL6���+��f ��֚��ob}3�����BB��;aX� �j2g=��B�҄��8\BB#fQ�HҎ{Zl2#������`����{࣑"#�X����`����~�Xb���!M�"���A�ؗ��::j�lTT��^0XPO��P�2�����~�_��A"���z{����.\�&ȯ���q�5E+�ӷJ&���@ǫ���]#ޛ!��ƅ3��z<����t_��:��О�\`�������S�E:���2�'�xx���{}=�w�:/9�@�y���+�,�0_kX��ɉwp*m�����36%����A
*��ȣ$Ez���K�򞌨����0�/͵���Fq}�_��,�[@Dt�^T�x?69��\�du*�!UR-b����x��e�ӕ�wvԌ����Q�O����o�)�"�H�X\R��%P���6wJ[>��dMD�;ЏGӘN���-9��} i�}곐���h7FD,��ǣ��?�(b�b�w���f�oiL��l�e��������9�����!t�S��*�')0�0 8����i� �c9�O��n�F�C��tk\Կ�bv�t��r�U�����9�n���ng�>Y����\�������@� x��$ޯ������Lc #��2�Hgb�h����X6�����@�	z��ό����nw�!vI��9�)k=�_����-��-�(�&o��+��4yrA�=O�^M`R���!��u�2�.�x�yJ�o�m�s���@���<��6P�@�����kf/�#��ߣ�4�9�D���+�^z��ѥ��� v˕%%%
}?t�;K�N��3�s s�O;�] $.|m��Qu�UPZ:lc#&�u�;�H���k?�$
��cԴ��#�m����=��W@� ��U,�sx�\����2;{D��Ä�Ö> �)�1���`��UgN �f�R��x{���~�M��޹��r��ʅT;g^u��n�N`$Tq]�n�/���[d}��i,�d��=5���1�qVTy|�T���_��y]�Z��}x���Y1��y���W��a(1�U���l�rpR��K��X�vp�)������m��1�'~�c�񤦯��-�F�C�Q�ٙ��@2B�8\�.F�r8ȫN� G��#�$��M�K<����=��rM�ߤ�9A����"�k<b�F�5���.)ybhh�{PT�3S��) ���v���9dvbC�-��F|���s2�k/͝�S�j�ÎD��ᦱ<�UB�:��h9�a��j<Y��x:�������)oh��|�Uggg�MB�k-�(ٕ���@`�.�r��|}}w��/dЪ��+�Ѵ��[{'�Q9cK.��o��uvVVk)�����7�B�ȈT��t����i�B�33���?���Bb�7�j�s�=XЎW��H�ha͒h,�?P���ֲ�6�24�C�)�ޑ����&���L�����M�Ƒ���5�W^��U���}Y`�S2t�LYw2�ё����R2�v�`g{����_�>>��Wth�����e�T�w�Bi��h��Vǧ�|�y��B�*g0���J�їn��h2w%sYfM����!}a}TP@�4�Xc�34=3����*8:=�;�nN����	�u��4��K�Ĵy��{PFJJ�ׯ���V���&6���
gS����r���[�j�`���pO��.�S,7Bs���!�[�%X��~�P��J�I�,��n��/ii��,�<��y}{zĺ���P}�r@
�������)���w��Z����������[
��םKGO���vi�_�h��j�<�l
��t�� O�9�I
��f�1,\�%�2!t�j�{.�U5){a`@_�~E��",z���������𘳯�Y �G]���0S�R�J�1*�o]��ݩ4/�%���[��q`C�8�T�2X#}${��t �c��?��pssgegSQ�����B	2+�x�jV]�c,r�����ݯ7�f5��ѻ;�"ޖ��
ӫ��_2��z����ƭ^�KC�y�%�"�6��ǩ����s����z0z_��P�8F���tL/�D�S��|��MUC#�")#��R�%�|�]�H//���Y���7��$�]tkl����������qm�t+��h�SD�����%�uvu)]�K:;;C9��qޞT�9�\�B�����_�|��!x~'���G#������Z^~���M���,(���|�
�b]�P�׹�H�[xd`�#R1��\^�k�]�+���UQ��+�xK'G�n`�����⪁��]�԰�;r�#%%%9D[4��Ԑ���&��֒ ��Z�76���+�3Vl�vq�JXubZ��� ����5H�����Κ��H�	��l��3�Q��*)EO��:�-,(󠠠���Hdr�a���c�-����#��� ���Uv�9:r0>�+..���MJ�����+��ׯ���FG��|E����JF��$LM����E�jkkW���Ӻy�g�ܠ��<�ƪ���7��q\�DXbѝ�ﶹ �[[�_��dt��E&��/��͠��e� �&y�rѾ���"f�?q�7�&M���8�#uP�n� �E&=�5A$��j
7Y�����V
<���?0���sZ�%�?}�t����_�����C��54m�9!!��:�;s��4AT�ә�Ξ�ܦ�9k�l�pF��x������������ظ�A�(T���-�Z;b�ޟ?�PPE@��� �� t~-�B�:�s�]�b|�.6�OJ	����2��Zw���u��"�B�㵗-��xB�k(y�L999�����ά����0`o���G&��ΏKK�HVDNVkk�8==�:��?Em/Q�e>���rG�H��$m�y�_�9�]��r|����s��ҷ���ͽ=i'��443'�q(333P%��:3��~.�b����7
��������	��|�}�N��`:������<@ڞ9�Xl\]��,@
$��~l��J�uY��NAދ���j���6��A2n��s6���b��[��{�\+��gl3���TU��f���E�'&�l�TTd���:�^�$�Sz���_������>J{0h\�� 3O�XĊ�n��]7����(�P�O������J4!��x�t
_L��Tk0�(s\�A_�q��/&z�I	Q�z1f*Zn_0�>��(ς��å���}�};����e9��'�G _��6X�swu-C\���f���;�pw�;<6���+ُ�Gu�SS=�m��E�I����D���"#ш��C,AN�A���;�y�#�ƞ2�~�|�~�T��r�!��>�EÒMʎTгD���\�����NrI��^II!v���2�[q��t1ODno�pC�����4V�E,_����i�'&B�9�ҕI]Q�����4�͛V�4��N��F94_!��A�
��y���:�	�iv��iZ-���̺Р#=���Y-��`�b;�LI7X�K��_���C.����(U��VQY��3(BO�m��8j���K�:v}���e,���1����ՠ(��&J-�����iY.}&���r�Q"�W6������[��f����_IC��{��=���w�W��-f�����=����K��n�����{���?C����	:��ɩ\G��Mu�:R1??t��E���g�z��3�\H1ç���/��Nl�4!�p�����dօ��
�&�[ ݵ��O~x�B��<���x���N�Z��u� ���Ԩ0 D```�.;�A�M���E�^U�����I��^;/l�P��pSdK�a�L=TF�J�	?���tpx��8��	��;Q[�������Q�\�M�O޵���PS�s_��yM-1�z6RQ�(B��>lQ��S��=1�/x�a��� Gˏ��̡)ޟ^�Fn�h�CW�Ʒ���z�>Z��E�i�ǻc8�2�a�'�bVi)���^�U��	pG�´�_���[�!�/3!X����::���N�KV4'(�HV�ZR"� P�`�Adt$:-.!a�ɦ.�m�$tB�i2t��\%H7���>�ؼ�?�QA'Ï���~�Ĺ/:0�>+[��-f�CT� �pZ9Czxo�9��v٣�˧65�/��'D���k����dG�p���Y�~�I<�
D��t��!ظ���e�[� �С����
�d���L�y=P�)������tYe�X��EA,M���������k���׊f��#�����#cc��琍e%���9��������k�n���F.! ��-%]�!p�)i���"��H�tK}s����u��sf�<1�g�I�����p5:U㖼��^��(��_�~�UM�]`���"�355���dė/*]�� ���O��aY^�]y5PYZ��hv���r�{-�O�N��襎����C��*ދ���
��,��K;����-Ye�����/G����r���鍓��zAJC#�f�J��
�;g�I��Ն��h˟���9��C*L���YB���kP@P�}�f8᧙��b�0RM��u����ʗ'@#��9(**���o	�WTp&�l�����}s�t�2VP�W�?k��yK��0��;�ؖ�ZQt���/�Wz�@,�r�}�B�_pIIQC�	wqE�eU��rφ�[�<<=C�ɡ�L�h�yн칳3O�{"BX�TH��Fz��P�D���
���_�`�7X���_��~�K�8�4MMI���X���U�H��4`?�8\!��	��(+�����51�����"1	I�:FI�<����l�>�� )�N6�.�\� �u�������ɫ��W��2��ߊ����P�W,��󱘚�w2z=�u�<��*�P�z51����B��{ ��9JN���ʺ�����5�e�d1���Z7n�UXK�� �!?�67�y	�f)T���	�2f+77u��>��Qr�>�P�` �{xE��4ld#��6�����z�����t{&�շ<�8k��R�͞����9`�ґ��'�b��`�� ?�-Y�s��U��,�o8�΋$@ђ�$���� �P���+���=�Bn4�V#��xef���l���F�Y�Ğ?y��JJ
*E��/�_��yd�J>(��%t����/���\�:Ɏ����1���H����� $�eq-��>H����r0+WX�����g���iY�)�d�eaa�O@���kH!�������n���f'(���� 'J�5�aT,
�UK+0�����Ӕ�j=�iZ��������BR����ٶ�m�i��S$��1*F̴E�@��=K��Ҳ]�EK��&�ҏ�kzc\a��;5��f��74ނaC`����Xn���zd>�?�T��H�"}->D-u�N�ʊIL\\�>��+����݌E`ވd�,,1����*u�7��.8?�@�Vt���e����^�.Yt��Ȝսi�%�H.b9�����.�?�DlllCccg��O�<	G�RaUK��X1茈���A}X�����p����}��*���O�G,;�Yh�'�m��Q�X2?�Z�V	Z�G�p�����\���E%�̌��<�߾��&����D� ��!Ζ�#�k� �@�8��Fj��%k5f �~.��� \�/������]Ͼ]O��*>�3Ʒ����k��OX����s�r�Lْe��ѣ��׶X��_^�Gٞ��&��G�>��:M.,���(�9w���	�!���a@��?0�o\�Ps�Yc���gt�.x{�����م�P����~8����@7��i�rdl,\�����6?�/��2@5�tuukz�o�m�=��a�cm�/eś���B:eA�BZ4333��-YI�~dÍ��!��L�;&..X�Y��P|)5��2$�I	@�
3tI�Ym�	k-`z��|��H^�E�}ySPR�=��d��������c����������c!h��b���'�B_T��䃝UE��+�R��z�|�ӝ���>%����7v^)nݷ�C{(�s��������dzI!��pIV<϶рӸ���ܝ��{ӭU�@Z��"N�h�f���I��$}�65uW�ʺ^��D��qM1�-�7o��v �'���阮�a��N{c���;�e�)c��w�(@�̼4�us�+�ܳ�I� 226nP	�#n�/�����V��Zss�O�Φp�a�z�4@�B2�Cr�n=�����jo�d�)V����0
��)*--,,��ZJDn$eif���ðw��RNE744��x_B{Ҩ|�����e����E[g秆���h�����P?�b>���J��(hS���<����Pa�$�IzI��D�}��������_�p�A z�''MiH�8sDD���0(�??�^NN�Q,>��uE=r�}??q���a���j��E��x���� &�p��&�ɛ�����[�B`񹸸� }��_#'v��ÇQ--"@-M�Q�}o�'�6rW^�W�P���n�/����^�n�w��`��9w�ųVk#�eÜ���+#
+W���W��Ϸa���o4�5���M�)A�:��gC.6W�KV���8�[H$Nk��\�.�K�Tj*r�Z��5�-*t�:���޸̂�$k���C] �5444#�t����_i!:�`+})%��i�Z�Z��T!x�VSx����f�V�����S_�0�[ܦ�:�??9ʨ������oMM�ݪ	�P|z�������8g��e砱����M�������q�K�}�Ny,��� �U)Ӟ�<���S�S��Q"æ��S��m�����r3��e��p趉�:B�&G�F�8���B��ErT9��{��4�U>��f���ݻw��$�kiK���,�ǒ���0����?;2՞2'�/u ����܆��h@�-�If�sf��U𥹹�����	 �x�F�s7����#�!aT�T	�k��PXK��&_�݂�K��k0Y�N�����0}R?P�)A��/E����^��W���	[Ђ��S�F�gŭ�QC�֖{�O��ô���;`a����͕-���蠖i����w�-)i��f�I����OB�ٍ:쩐���o٪62;��J�c���2�"驩�J����tttP��!��~�'A�et�g����Nq�6�|Lm]�<ݯ����J�rϹz�i�Ώ1���M��M|}*���S�"I�iד��ErЕDx`����S��� b�MO3p�Gs˺�����v�N<>xF/@�z�����
�+�#����x�&�_�=�E)�[����g,�sr0��ӆ-��$�x�6=}��D������W�bB��X�Cjhn�z�&S��R̃us]�0�������Q~� ��t��ϐ%tBt<E�;�tJQ7���4�$���������g쩚!���V9���.nn�Ϝ�`t�M)��d"��Ɯ�}�]�\��ED~����@7��>�p�\��E�����<Sr~A����e Ƥ�G�������홀��3����y`t�]u��K��S�r~�����rl؇���Ұ�WT4�V�]�^�$� �|��&<�X����l�Je�ς�=�ۂ��2^b9��e�EpGFFj�8�ْ`MdQru+gf�o7m�����%]�]��fZ�N�`c�hDF��7�c�U�0��L��_�=�z�;��v55��P�XS��+ί���Y�^�MHX�5���y�~���o�B����&��+�xZ=��)�>�T�� ��r��[�PgG�tt��o	˗�Ap��Ąe�du�^�}�{��x��T�
NN[����ksH��a���D�{=ލ����i[�p��A��'n�*V�vg5|�[���E`�L(�6Ws��}�76�U���wu�^�ZMfU/���u�_�9���������؍ F����tt-�Pĭ�h������
�"D՚���6x�3�o~�c����j�[c H�yXN�H���
��X���T�~���Q N���S�.���-� /v��F8�_Z��9���W��^�E��
?~����IӉ���|�̔�{$��.@�M�P:xi]�F���m`�>t�I��iE�.@��r.3�����/ے"Y��
��Wj

���n���&�1�î�s�e3Tpwxu�����WH���ʳ����/)))T�'-^�����dT��ײ��̛�kkj��[u�חp������~�AWOw��S����ZK�H�V<�c�jaq:6�����`V�%����fx\�|l�I���M�P��X�܄{1!���6�L�;9��"<wdn�x<S�C�v|�ܹ��,�j9Y���}1�>@���Еh��q�_����V��OL뇡��O>�7h��R�\����js�8�*�2�@�=
���@�_�!�YC��~.��Q!:k@l���+d���9	�/���UtBa�v�P̚�O� Q ��-X����qf�`�Ϗ�>�^>��ppšvd�Ǳ�����i�*�uI-`C����~���z����U �I�������Qa���{���W/�ii�8�A<�x��܁�P4����0X0��N�pǔ��攈(;�Ό�/Cg3��\�cQ���ڽOEN�	�j�ӟ�
���2ģ޻�u5-�~*�,LϜJvJܾ�O�#��e*k�
gft>Lg򫪨D��&��'��C ��d_V]�`@.��DCr�+������A}�M��l��������n*܈���7K	���~gz��Q E��prZl�(�������Hٙ����}P<�$Y����a�)疠�����-�k
�]�f*m_�Zq&��q�Ȼs{GxB����Ůg�[�w�BuV�@�)} q����'�
5N�ϡ������&���kZ���FzhN���i;�{��3�i�����h%[>�bH2���;z����h
�+�T�z�%�������#���I_b-���b�qG����o���,��N��TT�|t,~ݢz����;��Ö|�;�G�{�ZZ�����h�x���P��9uC���;�� ��fz���>�H������!V�p��<*��N͜CFvv��c��ķo)�-��_����}���Cu��y�ٙ�$���� �� �%�'��Z����>���]��ô���������缽��k&�ϊ̲:n�[!ʻ@�:��')���sp4³ֺ�;��{��X���uV�����l�Z�۳������A������*�x9b��=�YS�6���C����#�mƩp����_��?9I��N�0q�\=��@R
�/����z���t�Qs@Wn,:���1�<#��0}�������m�e2�����څ���\��9�z��4����7��A9Kfn��Br�ۅN6�;�Vcx
>~����:��=��S�P71�==PK���8j���e��KIF���LY�7�����p�ќ��x���i��ΞZ���ȠR�N��Q���F�t��L���j���Xx{�(j,�<h�����x*��F�9j���uL����J��k�x���#�l5�P��z�&��$���N��y�������e]�Q�X��ۇ��e�:�)��=o�D
]�r�s�˴1�= �$0���w��&�ޣ1�.�5��ۯ#<��5E��?6�˜��vu%P-�W$ؘ���L�|uy9�P�sR���#�1f�� �J�!��}�A��פ�:��Z�>����
8
�a��O��������<���V-]۟�}�VRR"�(Y�bY�\�b�����d�R�Z�<vg姙0�(JOK��a�]���~[\��z���з=��q�n!:9o�8���ׯh��D�M�8-�Z�?|x3���:*d���-�8�k���O�	��^��D�Cw�y��aY�4�WW���$+W��e%f�����Ee��ͺ������n�x������v9z��/���.#��׿��ĕ|L:~�㺏١KI�h,�IM�~�����mc���]3Kn�o�β���|y?Wy��f�,(������j-�e?`�jJ��r<����wa$���*s�`zg��TGECs�80���Q�=R*R��K)�ki�;z�o�M�/�Ԗ,NBB��GYB�������uW."�ڦr쩫+}J��kJ��ѣɥ���1B��3\�,���	ئ�G�@%� �{ޝ�t|ǘ>rxZ$Y�R��i>,R$���ߔrU\��F�1���i;����l����!��^�F��#�����#��h �����P\��a��ݳ�D'ѱ >0�VKKJ���<_��4\��N/V���wťǂ	�:Ⱦ��I�&q��u������σ�����|�fv'5t����� �RRO�������4>膳נ.�Vij�O��t5�z3��УR'�0C��yfjj����vK>};����M��Ö���C�Ԁ�KJ�:|��	`G,��N��9���;�R�u�-���y�M�_]2�v���S��Ӈ���(�<�f�T�b��J���?��H��D���Z�H��"��{�^'���fh��8�t?�����3���/�	Xd�t�_��B��۾���A��dKAh�D��&j`hXtH)�����PCW�猋�55o�qE��S�Vg%&��P�yC��]�����~����Jn`� �x��X̬�3ml|�A��DS5l��-L���o�7�}��' ����i�Lf��utҎ=c�X98�E�W^|�i).f
|0�����^��*��kER�|z���� t�/z�"n�l������?�0�΅�r���i�(���;\E���Ŏ�#�l���M�l���#��·+4 �]DR��>_�:f��[��
�Y�"q��ޝnHxV�7��&��a�z�=sC�~�{c�)"?�8��<���v����q{'�p�� DDD��V�
���N*...��<v�ɹ9�j ���=�5zV�OZ_r�:Z�&*Z.ޛ��5�yțf������ �I8���x<<r�$PD�c��]����]�����3��o'(���TT���w/�uK�+�[h*su�ć�&K�(��0���|0{C��i�E���8T���������tS}�:�ď��3�*��q=<<�F�v`�)$/�=G1ɘJ��{��8l�l0W�6�{���~������&�(��ҙW���z�� QNq�ш��Z��U�}��$�����E�˪u�Td�}������.i��q���������3����_��'c��$y�#�Ҟ����ͤ:b�b�j��P�� �_��;|���#�����6D�鯬�K�D���O���L��]�M�F���Y�������CA?�̴ײ����KN�!����hV�?$�z��FUpXu��! ���$E�e�}� 	A&�W�[6��(�!I:�i�sb�w��_p}2��@u잙����� 2¿J)��k;m��\�~-U#s<�'�_�����3��	:����������r�W����l��~9?+�j���(d��X?�]�(�S�o΋-�(/L�J#�Pa�s抑l(mEǋ]�w^3}@��J�G�}L�O;�Ah -Qi؜t�
�t%f�r1a�z���KhUa��C���:ւj���&ў�!��6:]�??����:昡c5���T�h��9	��.�'+L�x(nh��Ҝ�E�:�o)	���ekʒ�l$$� p���R����������pc��E��w-D�k1⎍�E�ʁ���[�w��}�,�3�eX��A������Q'�2&�&���iw�Q�@
|g�K[[�I���Tz�Z>>cbbؖ��gz���I�;�����òÝ��ɬ,Yb�5�T��6�'�#�r��o���b�mf��AԖ�܌�|bq1 ח�1���ܴ�G���[:����(Q�+�{;�Q׉��Rl�B�߾}cl̰ G%�y �v�ݐE'���B[gԤZ(����5UY��B�=p�'i�
���M�xf^���߯�E�h��9>F��ϟ���٪,i���c�-׺�nx�M/qN�Hn/:��X��MJ?_�%�o��͂.M���X^ ��K608�va�v$����>�>K��#�4,,,Q2:�;h�qpp�����Ġ��d���~%��+Q�"����h������IH��c����Z�H �d׈��^��A�,��Z����s=V��O��4#u���w1V�������/#ؔ���o+f��e
'ѩ(�|�44���33�A$x�<��Z*���˩�b��I��3a�S3��G�|Y6��y�V��2�e�y#j��VA;�݉���Z����o�E3��]]��{����C���KC$�t�v�AD)x�Z���łQԫ�Qdl>��j	?���J��0I�9=���L`�\�"��ȴ�H�/lЕ��sLI�%���/�2c��-�Ik�8��ٓ��^�b۵�/�DAf�/UC�����Ęϗ�m]��)�����ry�{6@�A7*]��@}ɑ_���z�4R�bn�����^f��ѡ��|i�L[��i�;^�xArr���~��V�~�v�9�?������uJ�bؐ��T�ޞ���k}�K5#��쮇iv7�Q�٠z�������%V�UA�D�듻%EE�zzzB��q#.�g�83U�Ա�_SZ^E�V���Sp�����?1�>uÝ�� ������V��}@i+�D�q���c]�qz}�sܞ��Z�mS��%�w��D�l��.d~gbgo)5���k�b؇8������-a����,Clu�D('�{V*���,�j��x�j)��!��ϵ��aЭ�`�F �r7�pC����������?F~ʀ��V�g�'u���?Y�qkw7L�|`y��<kM�ڕx�=$����q
"9c��S�ښ�O�,���2ZZD!=f?�IJ�n�����'�c ���3�������eK�	>��b�4������kE�:ߏ�sP����$�������Ch%u�V{�W����Bf~��l4�{��]�C�!B	,�#�4�NJ/����1��u,�W�?
��L��޿x<���gL`�����i)G�V�\]QA�/Q'f5��w�A^ �9��RW ��^�j�#�U�D�V�ׂ5��C�y0�D��{��4������Ъ�=��i�p�V��g���fٓ!~Iɜ�[�a^�P& ����R'JT�t������%B��;�'a�!��j��[��.��Z��~��s�\�r͗�."!ݷ;��frQ]Ŧu���iI�PBe���\�ɟ��,|��x�)PѤ��ĽaXd'�R���W���LL~&�m��v#��+avЈN.#@!F��ٝ���P�ڜ��Q�	 �I ����V1�QcY=�,�s��|��	s�{�%D||�����A�~aGGG	w{^�Oh�?E�!x�}}��9���0ɟו���kO}y!�&�� �&+{�}E6��|}-�ks���3V�;�\Ê�v �����[gth̈́�444��;�Q���nRM�qķ�������UAr�Ohy���ѷ���w�>{3`�!u���ݹY[�:]�$����a�Zr�u�y�D�w=N�?s�,ہճ�� �6q�YA��i��{m���Ǐ���,�8�3�w�$����\�j���,+Ø�%����T2Я}�B��#������GL�\�V�r��2��x��g��@���5�녲,K�Ŭl«������BYRHːebggo�����jd�pJ�۷��>���_aa�K�T�e���[O������� ��},����*\ =.�Ѕ�}��I3�M����s&�X�Ԕ��D���x��.�[���ѥk�\�=Q`;x�C��.K߮IG�p�!��R�D�k��� ��\Rg�����|UZy��zrr��P�Ls�+	�	!o�H�[�3������&�)0��E���OOO�g��{�N�����!W{�xH�RE��bb�Y�9Z�Iq#\�Մ2K�d˴C�D�fX�%jo�L�������8�\�d eB��,���	;-(����]={�EI�w;���#a'��l kR2��,�Sc���RBqi��t E�8/u�4���umy��������|۽�vR�'�y����t�''���;� bdk�˫���-b�i�{�Xf�+(�/����92�
n�z���Ag��BEEu�5��*z����1vh���ы�h����>7IkI0��@�,�|�j���-���A��T�YS��Ю\5h�����V���qj6�(�v�Yc�@AII8�H^��u�Է���!x�*Ic%;d�ux���������?�p�*�ɽ���5Y*�P�c����߯��r@T�I !-'�n%�b�Yki@477Cg%�ޤ�� TkeuM���2B��v�tv�$k%�9X���[�B!{��"���G<�㸷�b�x啹�x��8?����LKKk�=G�5��'�a�2��.���_ٹdQrЖfYY��q�SrS?𬭭��ۼ���. ��P"���0:�[t��Q_����j�WHH���.�?4��777Ho����>�z����F<��'�yL��}й����й+*K��ǩQ#х�l` V�=]����w�����


�RR���+T��@+$�~mus����/���P��*Z�(�6�����F�I����!+�@�����w3�e٠ە��?g�[���J�s}����u���-k�8(�@
��R���>�8;�lhj��^}^8	e9�ۨ�?6�4��G��Q��+4�J����s�����yE�=''��^�R���q�M���$���e����֧z3��''E������~��*[{{&^Q����DL[�.�o��7%���+�����<��6ߌg�둴��!+J�u%�kbD��[����	WdLRm)/�*���$=Z�	�[�h#-�du�Q��.�N�jD�q{��>:T7��[�A<{&{��;�AĤ���J:���qfmc�OEg�?�s�*g������DF5έ��ʨ�9(�E=�⥺�5��������1����]9ey߿߫�^̃`�&Ib��b<W�߭��\��g����vj~d3���=����l� ���]Y0�׀�^�0`�S ���y�[t,���3|0�����MܵD�n:�����-�2].Vb�|i�?��3�DZP�cŗi�! �q�Chs��f_&��\�Vg������d�V#Hpux�*N������;��xr�/K��Frgg付��Eȝ}��B]��6;���8?56�ጡs�h.��;AG��p�6"�b�N��y�"#��ͫ��޹\ʑ�/h�\����=�;��Ry<���;;b�*+���d����v�k8c��.5/��r�za��*��4��,��w>\mmH0��k~D?��<������ qy��>=���M��$�����w4����צ�h9�뮿~�d���@��BU-��Y�1WVbZ���g$�,�z,j�0T�������A����"B�ⱝ4�O ��gۄ�ȱ-|}�v�`�l̫��e���B�˰uߞV_��Q"�$�S�Z���0��-�_���C'��*>|xZ7�'� &�K,��N��s��z�kZG6z��K��!��.�>���n��!� �X*�D�GF��^���1�C�s����b_��5�c�&b�����Ku���i(���_.�'^�W_�-�8(H����=:�3�Wк�h0��U�ѻ�v��hit˺y�>v��! ��4�Ö��m�`n$��D���B���bƭnLo��q��߷��.��� 7�t/��%��*�h�`�kI�I���gj��H����*u�LsWM�P/�w��	�5׺�Y��5��XZ޼4�#�qbRa�:Z�;=�j�h�]�7���K�J�=�}�L=�G�r�ٔ�:�L����kj���#3^؉���iD�
)�Y85��M��
��yt��]	�u��˂9�n�پ��A� �S��2�:s}̄*'���D)��ۃ��y��*վ7Z�8���Y�gT/�Q�Sp0�6ġ=�����||�_X\��/�����i��X�L�`o�����K�5�~x�
����R��3���ggq�A��A�WTT|���n#E���$��M��>{=�w�9a�ZJ$����V���l5Λӳ� �ۭ쩘qqq�ʠ���4MN�t�R�<�|2ߘN�]M�9���v�_��mβ��EƐ��̢�y;�8���K %��W���M�y��t=��!bQ�uӡ���eE ����F�{Q	�����\?��ϡ�+]��c�ݏ�S��@��C��K; �����]��E �[�r%���3;N��Db��-����lM�c?������uVn�����,.~ہ/�z�K�ȃүlm�o�V����?�@����;�2%�]�7����P�����:{��G�xF�-����3�e���X	��+� ex�̧6R�UA����ļ�K�<ENLF�6A_j��Ŀ{G�Ņ�z6fnN�eq/��Q?�}����J/�	Yt䝳�f=��-Α����^�����B�w��%�����E�q.�(��;�]��,�e��>y�g �*���:4�`8�,jh>+�ߝ����ڑ��zi�*�Z�w�/+}p#^.�<�DcNT���sMTD�N�⚌�+� <q�k,(..��5�Aŧǝ�6Et\�q��=�o���cyV�:59=-�������=m-��/�kh�.R�d�
�^�ӎ�$�|�%Fꂖc_�Ȇ�R��~�������E'�i~Z8#d�<����xUۂ�y:O4u6/f��R�k�阘ɱ��3�32>=���q��0��f�釪�_���,��7������Ap4W754��`Z��v]>�G�#7�c�:�+��z�'J��rߊ�u��P'^������`����֦913�Q�G��c"���:�/E���%�gH��\�ұ���r��ʡ����ޞ�B+g?ά`8�ȱQ�L��g���icƯ�G�ᣣ,z�5ϛ7��k9q��>�����4<�𿫨����� 3����-�z��e�dnK57�r����p��M�[`��<��Qb��m�ʆE���@	��Ę=+.W_ Q���iR?H�L��[��N����-�`�!Sġ�w�=FNM=���O{z��߻On�:���||7�nM3��0��]RIH�8[�OD��%''����MX֚�Zg���i_(X���%�IE�!��"��@'J�]�cQ��1����+�'��Ȗ8��C63�% ���&X�࣡��`�J��1���i:���j`��Yֿ��n^���$��c��U�;#����㬞hX�r1F�j�=�Չ�����=��#���Kd%_��&���:��#���3g�70t{�c�=����9����L�_�ˇ�Oi�F�\��]�/���	{j_z�p�&y�T�������}��1�P�{)�����ԁ0��|��i��)�Ğ>�s�uo��m~�(�'eﲲ���3�Kb�A鹶�@�X�ɔO[E�]n����]?���PP�������/�~Z;4��D����������E��H[w:���Y{�|(>�(�JR0�z��Oh��ϯVίb(���Wl�<6��z `a�6%�8U��������Ķ�6��BB�ѫa�]ɸ���bZ\��'�Z:1��+]�g�#uM���gwHF1�aC�'
'Y��(��toe�Z��Ó�؞|��
�4�c�\�ʩ5w���@���m�A���?��T�\cP����v�\��Տu	r�����qc�ٴ9�'C�)�e��E�/��_����7ŗzl��3�g���/7ғ���¾�r{��3�������c���*.X��B����%� �Нk�����Cg�u�`�ն�(֯�����-�䖺��n���&H���S0�8��u�{q+���-������A���{��"}wL/�����Н�!m����s�j����.��5Bk؀NJ"�3�����/)S��\qk]vk�ih`�>����q9�3����_��t�Чubb���P^������I*����!h�b�����W�ʖ1���𠢢jq�P����n�V����!;�Ll�u1¤�F� w_X$*�}bŠ���E�걑nX@���(u57+��������>K��:h�2����,��'���V�Z�265��:�˴ш;<���s�&�j"K���K��aa��5�u��BW�6;x�*u��u�b�����޿]!�	�\��ɿ�)��)_9��}�i7�*�z��^���GLӋ^2LJ�C���*	RR�&&u0
�QM�c	N�Ύ��$���ń��O���|�UY��f>Y�".<�K�[���8��	�47d�Vs"'nW�W��,	ί�/���ȴu�������i
��ؘ����2-�����
9{{{��gVvv���?TW/�.8	W�t�C|Pd�i�8�����FA
��1{h�5?�*<�������\�x$���sw���b�Jsp,۾i;��Ǻg�H:P�[��Φ+eDk݁����~@��g5���lX�0Nt�诊������7=�5�ž_8���>��Gmn��7��cv���P�/�L��P�.w �9/L��i��.���^��p�ڇ�ʰi;�"o`��bܤ1=��}N�/==u��1�`zzz�z{����I7p1m-������@��Ǒ���1��i��Ɔ��/9p-�����e;y>�B˺�1�a�����ۍ���.//�W?�M`i�Q�����[I�TgO}�\�Ph�O��髟��=��E�{8���D�ߙ����X��p�O�hk�����O��;D<-��h��Q(l� NP�������E?`Y��G����B����8k�8�������V�^566*�?�;�z���o�}������� E�.h]�i�h����..5��|;��p)���GG��L˴���7�'c����n�ki%��O.ӭ*��rB���b�����U�����9�y�$�q+q�?��:��j�iV�����V
^����|F�G�)0�RKdL�B>�<<��r I��_=u��e%�<? �x���!���4^w!�'2|���hu�|��jƗy1wbƋ��П��V�BY\���|�J\�;	�ڽ�����q�?(ʒ�.�k�G�L��ǕŚ@J�A{��]N�6v�K��=R�;.[΢�K)����a %ب�M_�U|��ӿʑ�1ѯz���������{�ߎ� P�}d$� *����9/�� p����.����䌅��v�E�N��p���Y� 8�Ԍ�(($D��D�Zz��i�z)/� �F��R�Ƕf�=&�^�] 6��DQr�1!��pv�,�Q�r���T�8'A;·���<�@����t��ÖQ4�S�¦��l�#`�.6�BT��|7-G���?��j:���2 0���$��f�i�5ٰQ���g�p�<��~�Z"^J�X;�F�@!��HC�Ό�[�ߧSnfO}%�NXƼU�qJP/�>��vcr�VpN%L���������$�$*2n��'>�WR�)S���I��G�q���߄�Rq��aX��9T�?� E�c�ﾻ*u38$���%U��ܮH���ݓ6��B�{�1�Y�k�5Y��n��!pS�Kx��% �w/��A'��\�:7�ї��҉/*��T"d�h���מ�SSI5x� V5�1�ZGZG��2*Q� �8G�^L��n��z*��M�0GB�kߗ�*u�I���Ǉ�@������\�9/ܨ���Co���2�	�0{����&بP�!~~~���l�_��Ϻg{��B!�.����v��@����,S1n���3�F�1'W,����A`���˫y�
M ������<�	�Q�p�>��_�) (xx�J���ӳ$@���>�;��G�������u�֋�/�	v=�<��1�Vk�Pr"�ɛI#3Ú
��c��A��{3�TV��]}��b�2�^`�`�^w:�S�!�Ȁ�b[ػw�*��%�����ұk��119�xv��aݳ�o��1����謔���u���td�ͮ3Tݴa� �W^Y�\q�;������j?/�i1i����.�ߘ���C��C��M/��e��FBe�%�]��wwK��;P<׋�vL4�;-�Z螜�LNN���Zuٚ�O�'2�&�2j��RǠ˒��+tԋųl#}�?YE3�*�"g��J���0��\w��d�QE�4�3-�<���㽎���� ���1��үQD,��I^�xD���7ww�����`����+�����y�Ǘ�� F��3G���&R����'�����<�����#}=�'jj	�)(ʱ����=�s�����~�8��/����`�,�����߿^������uN@�@z���������ަ��>L%�GɅ���H�a����=?&���� �Z
��A��M7���5$�"���M3�c�7�K�����Xճ#w׫w�������g�C9A�S9223�+q��)����e�SKvXy���y�R���X���Տu/�t�I��Nv�)7��w�5�ET6OLMi�߭�{���ق�@�^� ��z��n�Clˣ-v�j����D�Au�L���6TՒ!A�w�v�'08�&Pd���ԟ������z"e��W��������WH�+!��<0RS������#��T�Jl>���\�7�y�b\DH��(k2��R������\Y�p�,}��Xчp~1q��`���r*2܈Kz��;�?�[p����-C*�U����F�ѣ� ��,B}���]E����W6�����W8��:����˙V�U~�qz�CW$���8�R��p�A���F[3'��{xyAg()t��N#+�l�n�i�y�:	V�H\�?3�%�_X�tʲ��K��P��D�H��T���GX���zb���?A�|4ԋ��gh������ʆz�����R�V��;1:��E}�����c�L��{qR����@�o(71�7$]g_0>h�I\T-^��2�����NU��˺�˄�>��X��ve؊} vk��ս��v���׃���v�^������H����2��t���Idxz�+˙���V�إL��#�9�+b@0�&m���Y2�����õ������"Ͳ��e���/kɻ�%��|||F����;M g�Zg��Ć����bP� �������Օ 7�g{纎��ɉ�h�W[�ZPPu!=|�Ӗ �<�j7�;1�8fƵëU�+0�@ �A�������&����,B����A��bT@`��Z�����
���<G�5�ji�]�k�Te�XI	si���b���o���;���>_�|���X�P>-!�H��Z:0 @�� t�n�V�4�I_�_��HveH��"< �e.ff��2y�31�˗ek���"#�]�ܸٛ� ~�V��O�Bg'�.n5oX/-L�}����P�2+��44d���_����y���McR-��]�p1h�B�Q@@ /9����� 5zC!���W��iS�s��&ݠ�`2�3�Y�5��Rg�����yp��>x��It�; }`�^�i���< D	��>:JMG6P$y���s��@q�CV�ʖ~�6�,�*��!��|� ��Ə����R�刧�r�����V�M�_#8�!����:N���s���T��N�%O��I�r[����뀧�{���ȖDF�&;������{��%E�B�ɼdeuɸ��[�w������^^�zq���<���>�9��ያ(���9����	bv�����.���Y��ƴ���I�?ƨq����ˊR�,!�}ư���ntH���j��l�ЀO%o�|w��r��ࡊ�
�z P��
��%�r***3�TyU��X�$kR���d6o��pQA���.eP�]VvrϞ�B"�VUz����b�e{t���-̟,ݧd\LJƖL^�;��P�n��	\�;�S�	���_N?� kK�d���nãM�����*|4򶶶�k��J�H��n��DI��j�<i˻��UE�����{�\;'�'���۵KF<�S�8�U4�D4{�}um�_Z�����(oll��M�]RR�u���cecÙ��I��a�PV(ʬ��N	8a-_���`���Ι\1<�8��DO�#?I6�d�cMP�Y�|�Z��_v������ �����"`��
��w�[3�B�w���?���Zy%#��Ձ�m�}S��p	6��^������-�\*��e��W���~*��>��o3���?M���m �-3队��ɛ���c̓�����ۺ������'�\E{|��ŤC�<��`x]�Z�8�:�w�_>*<C��D�1l���dffC�f������!o��@�	�9C�=a���~��v��~��Nxa-����R��"�DU��-��X�Ȏ?�ݚB���CB[�f66���,d- t������������ä��3=0𜈄�P@l���۾� �]�())�'�g�e���+*F���ץ��-���gw�*�H-�|��8�{�oi ���m�h��M��:�3�o�pK�HS�7:��|BB �fU���BV�@�P�p�cT���z+$ �5���^O&ϔ �����|���&��R��n�I}���3T��b���k�2ψ��8FOLL�~k����`@�V��ŎS����p�W�ӳp�@'E@�M�*Zjl[PPPl�y�1-/{ls H��co"b�V�J4��+����Qr�?�7��Ӊ��#E��-}Quub�^^�Y�3g��i��F�Mm��J\zE�0Ktbcb�Ok��t�k�xJ�'�jV\V�����:�4�hċ��N�s���M1�EC��h��|��4ߗ4��:������Y���g�� ���r(��'��Ć����m1�]�`o�����E#��>�tĊ�[����ڀA D
�d�h=�`.H��+.��N���N�&w�ی>���LZ7�L�j�OW[��d]>�,Z���p~@�A�v�|С�Qj��������c�%�ۘ�o"i���㳭N'>|ll,�U�]⌯c�)~�ߍ���H$�R�L���ʀ�? ����c��_���zu�¿T�IV[�rp��@O�gW"[��\ӇƩ��M~I����W��>~�S���a32CZR2��"��Ġ����%+���m�u i�4��8�}�(J,}��C�°N*ᅟ[FǍ�O����*��%GwR��g�!����Px�T��C1[}*  �/*�����\��̗!;	J�)\k�쀑�Y%wG E�!9���2&&�
_ܵ�{H)��^�x���ː4�Z�p63�pF����S��CCG���.o��70`�l�71��u�?P��v|�Zv�r�v��p���f ��d���Ņ߮���fff�f�����-M�<ey������%a��� *���c!8ɺ�������W��&BW�%�OIMx�h���0�S�o����-��-��dM�4����p���t��I3�d�����| _���n�d}�9`G�S�Ȩ}y�%{ �~���/��?E�?A�1�Y<�L�����������Z
|TH��?*�V��*v������ӝVPk��&z�J����1ۮuF�1Cg,��U�N�_5B��a�W�OϮr#���
C��_e� �N�B�KD����Um�M�e��ck��)���悫hE��|�s��*	"^�2'���:%?�wH���H���3�ΐ��/�!�sgVzM�1w���6t���ʹ�P�sW��߿	�^a >ĉNQD��Bľ�Z%�W�G�kU��ځG�05���C�A� ����i�H;�M�l�0����C�]a�/\4����_���������P^� ���j�-9T.
!��J���?��e�.���z����5��
��|h	`�CR7�t>'��K�J�H�w2�Oؒ')�s%}����_��ڎ ��MMM'[|3QP������<Y��e}�rg	 �1�^-|Ipï��jf���F���6�%ե���c�[�[�{�9�`��Ƥ~���Qٜ��N�M��AUU�`��۠$��'���g��fvvx!��ؼ���ۂ:��P}ԗ�@;���$�F��;6�ݵsv��_a�����:���D��zM�C��\QW�T��s�Ez2�7���w��_>}ֶG���a���=Ӑ+��F���&ŹAnD����Z����(�ۻ(Q�ϒ�'*X���+ˋ[ޗt_w(��q��Ͳ�q<@���`(O=��w�僕��S�
�r=AP��G��,�z=�������3w++��^a(e��=(m���J0s܌C��E[�7�&*7<1ƛC����]wO(1���z�Q��X���\E�恢������<������h���F]�@-�N�;<P�g6�P�5��CE�ן���@�+��P�>����I����Ñ���Ҁ N�&�a������nWvΑ�sz���O��{�ePGf��9;99�w:����Cp��0�yĸ����J���G�^ӫ�,d���	hJ[[[U��o���CC.�����:Nx��#�6����OEi�Y�k?z8n�UU�`٤�w���C����Y>�?`W�����~� �c$��3D�v�>���\ʹ�E`�^[. �YZb�.�Rק��,R7��|P�G���qCՈ����1��S��[�7��HZx�<�ZN+m�]
���{�^����H��N��Ъ��j��6��W�ͪLU��Z}j�;������֞��Y�ė{�}�?~�}(���Çe�(Ct�U汹o���R��}뇟���&�)�C����X�Ǧb��w�:[*,*m���7�����Fh͘}��nYqoqn�����[���-O��_x{�iݭdg�m�c%�E��ҳga E�� #>�ֶ
,�K�)�?Gj�i���8��)`P���� *Т��;Vg��,G��M����=��;|am�p���N�L���,^����}�֥P4S!�U��"UP�Vw����d�����/SZ�PrI���=��uI"2K7�/7�mdO����.N�R�.YK����t�[��jc�{�H'�ڴ~{�S9>�I����pW���wxSK�m2^0�R�����/�y@�@����&�y��� ;��jj�������b��H���M��{
\T���ii@O�!�����986���f/�+++��z�Gc�$���\y�Dj���\WwMH�6�r�`MZ��lP���S��	����?B���+<;@LL��9r�G&�B��<��yk�wdd$�����M=��J�5��~�����<76602���Һwс���*R�3H�i^K���O��7���g��}����	�+>11,2���i���j�g!�K\�md�r.���}����?���,0�}es'�#/��k�$n�U�3��QN�e��IQ{�'}|� �9�+�-�c;��v��/�)2�j�2$6�fv9
/�G�C톨�s����t��Γ��L���cy���e2=��F���4<�t� z\T �>��$�}��a�X�|B��c%�K���0�k���������{�j����\\o��#b�?���T ��q�Xۢ��xSX�B�scY.vv�'O"����7"�766D��h.�G��P�a-��O8����m�>.�����iii@��Wp6�캙�sOb��&r�&(i�xA�^t�tX�|ǲ\�O@�uO�
F�s���4�z�M�^�v_	�w����Pў%�4�)�TK�>���$�Y?���Z�>47bZ`�!a��zr_�b���DzNO;���=״��=�����8E�e��P=�[��-,��SoG��1&(������#����/.n���#޷o��&�~~~P9��u��N�EA�hi)O3���<��켼'u��\������;�=@Z�j3��{8���{�gM�ڵlQ���9�<|
�VQk�~����o1���_ėu�� ��E��aqT�}���i�eGh<�E/�E�7�r|�g�ONj��hc�d�N������1��N�rr 6�BKS�ݹ�l���7느��B&-u#���4��w��ئ�Es��o�^�I����B�|[!19y�m�N��s�c~�W9�p�G&n�[��� &����<��M9�v���oO���\�s��`D�Zȴ@+���3���ӵ�P�٪G~/-#:���IC���dA����``@��.h����P�IIX{��w՜EbM�W1�c�VV���;�
�/> �Cԗ��6���KY//!�L#�o(U��q<..hV3�'����o��[��`�)���	"Z2��F<��k�c�¸�F\T�@zL�uTpiq|D��gYæ�����8ێ-K���,��0�RX����
��:����u�������VN��\�p(�)kk˖ᷚBg�r�������獫S�eH{Nr4�6S���;=�����t��OLN� _p.��a˄OO��{�n?UV�����`�Y,)#�����̇_PpY;��?�	�����o����z+�G��ɩ�����M���K���UD�����d�)������[��x�?�J�4<6)��� rz=;(u{��??L]h_B��L�9A�&Q	
	)��[e��W��nS���q/T�e���Y_�਱o�;�Q(FG�����U�r��Cu0
''n�8�	��Q懇�fVV�.��|D�/^<��|���[�8�"Dxxx<����~?	���
�t�j���"]�}`y�.��A�Nlt4�(1@= c_�� ��{���@/��:O�۷��x���X` 6�wuu�"����=��j�SA�(�뗯��b���|Cs���Bn�Y)��=k�Rőy1�>AA
-��p���~
2���
���y����Ƹ,""c�#�f������ͤOS7��	B,�>�m��.!++��~�y��Ox�� {�S�ih�4���ʏ4��N��ΩQ^��*J�k��C^?d�Jr����6���U�{���x���
��m����mz���D)�6�����8���9a\�M�Iٚ�99y�Ӕ0t k_=i��H��t��:�����ibvlGk��}I�{@eCi���P��:���3([��L��SY�Ϻ�Å��7�;{�����tL[�T`Y��O���q'''%v��+��R����7�2��rC�{+��2������������[�K��;#�Je�[��������ݎ*�7)�m���K��m�d8A-���	�� -c6q�5fF�*CC�a���-�$%@�L�:ls�ɰ�f1�ej$V�k���L&�#""�W�q���C��xD�kj,@Ȱ���tfH��v`����Λo��0�hx Zi;f2�����R����i(�2���-zV�Ηɜ3�P���-����5�jޫ�:����ۍ��ǰ,�p�G�Į���Q�w��$�T��hl�FF۞�j�]]���02�����Ƕ(�:��]��#je�� ���/҈���d޻�_J�8]-���)�	~?��g=���b���j�R��lPs��lK/�"�J��^^^P@#`��������ւ�rR�Ҏ��2��Z�A��1/���s�/�1�!y������]�g�bǮF��v-�o7�����&|��(��=��xgG��G�&�W�;v���%ϻ��é�����A'��s~k�������)�d�������n���*Gff�Z���s��W�.�&0+Bլs5�댈STV�<�ͅS���w&O]a����	3�\����`B�
.C�HH�r5q�V��?2��/�q�XT�����l�Z����?�7�J
�Y���.9��K�X^f�a�Jxcjbhxw8uh�=Z�c!�	�uW���x���C�'�_5�K��4�W�RgV&%�-��]f�nO!���X������ӡ����{f?E������Y~�J�Ė�l��z�B9:6��+h�0іێ�~wڷ��H��`����K�(�9h�GӠ3�2��*"���]_�a�w���8����;�|*�s,���[�=�㧍�����pt�G}����/^�9�+u�3.P`\UKZ�x<���りwf�\�m�5K篽�g�vC��]NP��f3:���>Ȅ�uk�������/v���E 6/�O�.1��ȡ�����O�?�_A�'E�P��R�[�\�����^����'$��fd4���l��a��3�Q���IU�R�tz��ۀ�N����c�4��
��9c��,dY��.{��~�)�e�}����3<��ke���_���ᾤxQ*݇;d�غ&~J��%N�=��7�˴8�}�w���u��NӖ�d�wO�Z�%����V��v	i���|-�,s�g	b6Ƹ�{��~'��F��Jv��X\B��Yf%�B�ΥQOY��?*C]���R^W�:	��R��ѧ]v���@�E������`��O������v��X���/��Ѿϯ.��gַ���<����g�Z�ڽ/[����`��߇����kh	�W ������������?�b�$���y���Ї����p�'����k647���.��n�خ��hI�B[��!�}�X4R����Ç��.������8E� �|���T��4.�>�
P8����S�0���׿~���	�r�� �Be7���x{���khh���Ƨ��@�����
�1�t�o;xRSV���	��"Y^�"���P�ָ�"�Z�]c&\\�搱110g!������?��@�҇\�� PC����@��}fVɬ�������A4h�������lu�<Vd�������Th��������ğKH�8�����{�6$�@(<�u�	l���8T���	f�h��ż��aT�U���qpl{���_����c�'"f�9G��s1a6^�f�9��BS�u7UUuuV}�cX΁* �C�T��\���u��im�	
+8ux����^Y�6-�����Թ[wRn�>t��O�Y�L�K���8�麪���x�*����|�Q�k^WW�o_��l]O�(��B�8���#e�^n�Ø��n��-��� �w&�L����i�ZJ�r���h�%}�R��<�.������Ղ�о���X
U4�Ѧ/pg:$5	>��8�<=	��_��1Bw���KK��8��(,*
ډ�&N"}ٿ�c�x�iJ�)�	�z6�fc��e�gPTXxy3�
��tΆ�g�2�8�S�����ܺ;�������A�o~���`���$wG�{GU�c��9��j��KAZ`|���nw���k�J��������ڲ�7���kX׀�y<�	�l}��қ¿5 ؊9�wY�g*1���}�}LG���f�����R�ޯ}S*o(z����S4s�|�,����D�0y־���1�� �q�e%P�?�	���=�I�ǌ��a�t��MW@�}%jܖ���ǚ�qS�%=�g55<Lq����<6�kj���WQQ�-6T[)W�����l�vl�ڀ�����#��-u q��A
&�@�J@���tx�k�Cg���A���~����>11!)�f�ѻ�*AV��[�N�wUX����el�_@`�\Y�<���)�N����3����G�}�AF<�Q�;����+y1���LP��f�b�}5��ȇ�A��7�4�
��'��F���^����N�> X�vqW-]�r��](�lb���i�Y�y����oY�{����>I���`�c@6�F���a���z�S���O�Nfߊ{˿����z4L7Y��E�H��z�Rs9�4�뛛m���B"ͫ3�o�Ն�����gz�z�[xa�z� ���E��&(o�6T~������tk(c�$	�G��\�����������FF<Ӏw
@p�c&9�j�8�y�@���Iu%���7<��葲��5z7S�~����A�uL��-��޼l�Y��qm��j�����lÚG\"�� Hggg�q��>zeb�����n��| kT�+�,f ���"%��+�R��3\��?]���b1YY�@����פ��!���J������v}�����a���]��s����*]	������q�u7����G ��+��l�f�r9�L���Oɏ|+**��TB-�|�ԍ;��~��G@�i�:��Н^��MP�SۘC96&�6�;�i�͆.�B�Kj�Rq����=��1�XqC��Z��h���w2�1���?�$yC�Ws��A�f?C�f��s?���U��a�d7�w괹y��`7k����!\��L8��l������g��)*�@�/���W��r�)�A�I�ξǩ		�4D71�uJ����j���zM�us]8��n�	�Rޓ+<~/&��d�$`[�WR�V�rs�վ�2���i��bgi�J:�Ѽ�}�uľq'Q�EIE�ȏ���"���OA�kqoT�$�dt�&\�wo��'=<�x���w�d��-\RE������E(����
������^tDJ�$�C�oP֪�񮈥��(��v Vяʴ�\�L�w�8޼ ���:K�(k��L�6�X�O�����"`�0�My�|@�iii/w&�о�����t�������P��Iq1m����o�C;�����?o��nØ�ynB9�@� �u�q��П�a�-��瓻BM���q�-���#��R��*�ʏ%�ܻ��̹��|�B�O�=�Ul�=�H���sH��#���qiii�N�$ǌg	�� Ul_�<#�i% ���)4�N,.Z�1�h-3���
����Y��	����N���/!�j�L���)|�}t(f�1A�I�D����PYw��Ǿ����� �ޢz����S���u�"t�r���q�X�F����3}==���)�	���X���ѩ�����"E�j�D0�Q�js���<+��V�u�~�2#���x��"���[�聿_�U�obH�|c��sc�_@����
��(��Y��%2���[�u;
��� ���4�����E��G8�<��	�p�^���S{�4�4�碂W�4��z��>�Ot#Z^`��}*82.���ɶ����K[��ۀ�d��Ц�Dݞ�&���Y�ʦ�����)i�wyI���sch��Qn���_�뇕m;�nW��^\R��[D���7/�4���	i�x����/,,�� m����rA=���-�R���o^#���J�Xx!S->jd�����))]8S��)]q��-*㉂B�.� ��B`o*�]�k���(o�{��}���Hg'�Z��>5uu$�嫞��z\TԬ�1�A��<P˯���C�C�6�-X�V�M%�r��������<���IP2T��9X��E(���y@W]]}�U��iL*�������V�U�*�% j''�k4<[�Y�	}�+d�K��c�?ZϠ_��|u�G��7μ]1�lgq��;zI�;kY��n�qc�8��(�"-=��댠S�9V2��>"F"�w��鮆��~��)���s�ۯ��===]��F'.|����M ��A�,���!��9�---������������A:<�k����[��9��rN=��H2����o���6�L	k-��ݠom�m��]XR�:?�F��m%��%-�%w`j�a�uֈ�xc�V!�?�˪�-3�uMM�ö�m�����%�t�Aɻ=<�5N��&�ۺEkΈ��u2v�d%�������r���U��]U����ؾ����&1E�?����?(?�� ��9�������B�^4�[�kb�|�6��e�}{@5\O�·���'],���ۼ�w��5�8�f���jW���XP�� �PLdr�u��B�*1!��!dz3�~��Ն�T�cy�%�]�ӛ��[[����]��fi�H��W�-$�C�~VΥ?U2��E��(��P-��Y	ܑg"����r������0n�$��B�%W�����T&	b
PR�ʉ����@"�ZgwX��XƂ..�����ikks�vw'�u�V%�ʿ=�޴
�/�cF}�M���X���)�A*�~H��,�{���YZo�	U��ׁ��ԧ����?s�������rl��c![�[�8г�eg�	������צ����	�:W�"ɀ|�۰�&��w�i�7�0H����@�]�7u�l~@YY444{,ۜ�6�w�]5�)<<L���05L�& ���l�������u��9�&y��(@6��bD{T )�HV��n'@���0ܹm�OeG�n{Cɛ������rs���-�ڷ+J�:�V�tmx*|ew�4'����N�ɽcrX6�L��/����� m�w8��;�hr�b�M�?#��%�"��V�r��> !_����tkILX8
�Re�.sR�F��$w����R[���Y�変��z���^3��L/H��a�6��Y�#�E��U� �3��3jo9G�ɡ8K0?Q����x���{o��0��zIQQ�JWOO
`x�%����Kٱ<�S�A��Q7����YBe��X[[�\[?:�=�G�*��]'�ƾ+��g�g��!p�
��55눡4�\xEX��k�g��C]E�_wK���9˝����e3�{&�5fii�y!��}����Y�/AMI��sԌ3|Ϯ3����R���[��Mh�h~!�A��ܼ8�l�Ǐ{��O.Źm�_�ξ���xM=ō�&�U�n��גּs�H(����O�>������
X�a�'��"jsM	�����G������F�>@p77tCQ/����J��Sc�ϰX�����X���456�t�m?���������2�9�j%%QM��98�N//�x�LGC�H$�d�6�C*ݹ�h4_����wh���~�L��*�Hz�W[��6z��xkb�cN:���d7S�F�w��6�ff������TSW��^>tO�������h/+��c+���Y�]��4�
�Odc;, װ��2;�3���!Џ�n�>�=(���Ⱦ &�j	]�w�����"�N޶d� J�ym�����Ĥ�}*�su|��R!7���x}�%#�}xJ@JSӮ~Fշ�Bz�m#�v�W��%��� r�c��#�O|�A�!f���>/�����|q�	�yxddʃ�:��2@�L
�<�H�އv�����٥Ζ�Zߍ"�G���Q����؝�Hs�`��iޛ�����A�<��+����7��st[�|W�W.>��� �5^�_�!��j�����1-���ۥ�TY��uG�V�������uXj�f��A�VV�m��������͛7G�8|VG�K������Q�A㡾(헐��so�7�i_�#�z����Ɠ'O��գ�����*���e#K@�L����6]@r ;^��]�A�r�{��Ԗ��5�Y�'`��P���k}�K��>��K�.�J�4��צN��blgoo�Fm(a����(B�x&�����1~]Դ8s���D�A_�3UU�p8�?n,��jR}�����w3���/D{k��K����@��]܈2dd�p"[�R��*(�~���j����Pή3>8�ژ��k�B��9�k�u��5�ޭ�*���\dֱ<������	���_tO-#���s�Օ=_^�*���|<�l~�qxX2\b:�v�,���-�Q��Q@�� �	�N�Oy�g�9�B{��,��f2At	0�uK���'$&�����=}�t��N%�o{��R�4vyMM�����	J�k+++Y997�bp,����4*��x��0�� 'ww`9�5n/Jv�e���H���R�ک�  ��rB"oޝ��,��7y67%i��V6N�G�]LȿD������`q.D/.��}G�~&B�ԥ#
��R���+�G�-3��\��H�"������m3i�ig����_��|;�!�c�v��E'����h_��_�ť�*�|�R�X�Ku����^ɬ����('55b�G��n:˦�c�xU
�1����`��o߾�$��cA=��m�����ض����P9��?Oнm��ʙUNB.e}��Y�
��=ܰ���s��jppp��]�ϼ����4�[�-�x�q;��v흗����a)��Sv��o�x@8�o|m�>BI,ypU�kgrq��)�Ǌ�@�>��si�&�eݾs�N���05�w�������Q4BCO�΀c�g��������*S�ܜQ��ۨ��;�Ʒ
�ɯ������I	��R|�|�xdX�� ��O�=#����3=V"#�8m�n���-���adlYZ�H�6���q�&V�9�6����}(c
c�a�P\Rr��g���`�PgF\�-BކС<uE_�̩:�Ҧ�?����<������I�S��  �Z\��Od>>��Qp�wUݱ(D� ��ۋ���7׉��	Q�p+�$��+�*��o+�ݺM�lll$�=��� NPj�!����OJm��S��Ւ��n��M�����eKfL���=	x�����)Cdddk�	L�*_��T�PP)w�ˍC���t���|�,x�}�
�?��"-O�gb�[��ֻ�����R���Չ��F
��V&C��r�+-cX`�l7�>uj�S@�Y�VoUFQ1J�pڄ��ŝ1����
��pZ�y��ׯ��;��4*��&n�8�C�G���j�4��],�������I6�ލ�mz#2w�1�z��H8S2w��up�ƭ�v:��@_R�^�e@*����&��>44�6a��b'�O�!J�_: �J$��/D��wW�ފ��( (O�>;{�	��%��ĮڿP��ϟi�Y�������`X�Ӥ����Au:�OHU�b��L�


�w;7<��z��?�Lr��	��ܫ8�&��f�nt32�44��:솉N�8�	���*��G)��n#�近�t&0�z����6c',���\L�=)������ �j=� �����TUQ �3(���%��_noo��q ��^'�|� ���x�,R!g�\p�b�j�|nv�<N�RlWs7��@2������@=�/���p�f����Kdfu���J������ʪA�m[��˄禰������f�~���\.�)����!H�g�r��>.V��+)��|��g�S�Ϻ�l=���f~P>�	~P��U�J�e���t�-�ݟ�/�{P^��:���������R��W��-�h��2�����O��>u��<'S7P�4� �9��8��TTT�\��I�',dY���rDo�����46�p>{ <�z�m�%W���i��s!��c�n��%�WDm�}O��Z��svjiۘ�\{�>�5qᐳ�J=��5'-N��hW�%X#Tm���o��RQ����:	�q��immEb׏�oWT�G���6�n/�� y�����`,�^��$n�H�0�K�muu�����-���Xs��<�WaŶ�6��}C�A-U$�<��-�D�Af2�N�tPv�����˅{����K��$%�5�3���+��L�IO<q���!0�v��*	گ��x��~�1��f�������?�ڍN5�?�����pm0���8MI`�g׿�[4򇴡=F��,X���ʄ�4���@ ��q��<�����
%C_F�
� ����k_[o�+��n�Du��mj�C-���+D��~�1�F����/��A���ڋ�S��װ�g�t�H7'+�q׽� ���GuF�������QdL뽝�G4ccb���H"�*܊��H�;na�ޅ�,:�z����Ɵ�n/�Ls���BK��|�8H�O�㥟�)W7tZ��LX�	`��޾��ڴG���o� jj���.�1`�����x��������k��b-*f��RiоP+�i0Z�k�:#����\� |��[�ÖX>�ţIς^�3��&ֶUp_m���^B2K�
����1@ȵ�)##����i.#��o�1m�k��r���~y��j(��tlΕy��$ �!�%*�t3�Ž��OY������k?���w������n^������K]��7�0t;;< 9��U�())A\&9�`ʟ��߾ڨ\rv��17�����R�����>�p���oPV�IX�S� ǀ���K��)�%������+Mww��E��6i��F��iO:P����:e&�3ɩ����� �a�����j.\� �`Ȣ��8_^T3kxl��
�8�Z����\������\E�u�2n����߉�?��"p,���Ë��s�&�DXX�?��e�"�ЬʠD���n����n�J�ʪ��ꃮ/����R�n&JA'(�����n<}�q�b��ؑ�Մ����gޡ��7��R{׷�;~���4@�S�X<d��m�/v�W�����ᓓ�A�#�B@�7�
����wS��W�˶.��W��.π�Jȋ�U<`���.����<U�K�_�7D,K�xƅ{���,)�ZF���߽#�#�0��	�=\������L����?*c@�����ʧ�EO��,�]*S`����������AI@3�+������Q*�Mn*B�{�ዋV��rL	?��۬��^]]��Su5l�"<��Lxt4~�ȟڲZu�,
�TS8�B���������{	�>����sI��D���ȕ��ݿ� �>����'���L�o	@���4���;���T�"�<���;�\��a��+֯�����75O�������zM�cT~�칞�h�#~T�+0+���3�>���/�%���%���`���ɉ��gx����h��'�>�(�3���@z�f�O��8�b�kk��%w�He��;wZ8:�:Rz�����8j'(�{�q<��낭X�H@��	�������F�aZ슆�&����ToQk9߿�|�ä���]9K˜9��i��Ix|������¯����=���I<	�jTMM�w�D�_�ͧ�;�����x)������J�L:

	A{���������ڟ�ݼa`h�id�q�Hӧ�:�@K��������_Q�Ga�\2�������Zyǫ��GE���}�"�%}{B���0@�����W/��H�2���l,�oy�5!��v��{�NAEuSbu�%�v%ɰ5�)A)�`��JʹR��7�_7^���
�߳��e���G=�9�(��YNT�0̠{w�^�������A[���H ���

g74L[R~��'"&v�t��{yrG�U��o��2�E�I�m�/��&*���f���q.m�k�� ��''aM|�M*����h0��ѣ����%ؐ���i%Ќ�%�It��r��G���������Z&�w�{Ϸ�H�]̇U�k��9���Wf[��t���k$W�9� -��G��aJFw������4䕕	N�t��x4hsP�p?���*v���OX�j���Arw�7U��"?fz�e����PA~��"�֑\Ј^�K���<kKAM큸u�x�U�� �f�Om��b�>�c,/�"��)~�Fc-���( (�qF���ݎ�WRQ���a% $�j�Ɛ��<�\]X�"���ۿW{!WR�أ7�L�8��gA�Y1V���%M?fv>�Hf�i�ُp g�.�␬���$pn`gg�ҖQD1f)*�@'�/\|>�����_�x�h�˕1��ѣG;1s�0)�����!�p:F2�mJb��EA�g�$�`����a��>ЉQmp��@�ល���cKKKR�[)eYYY��J�HHw��06���a@�՚�� ^���e���Ϙ �Ҭڠ��P_h?E<��TWW�\'�}Z���NVV,˻�\ݭv��t()���C
-m��hr�0����O���.�;�Z���jJ��pW�t7��1���؍�/��]���N;x���[#o݅�#�N�Y@�.,*��$"c3	R)c�C�e"o�<zerC��}�<S�k�O2���z���s;Ĕ\!�Í7��`Y�ww�gw�S;,^)���J�w�,��E�$���='(���%�Z���kw�-$?���3���bs|�h4���\T���N��"�7�H9�ɴ"ϾC4�js}��9��@�m�ҳE�r���+���:��=}@˵}SfI�y^�,���k��p�]i[�Ĥ/X�*������J�ѵܯ_}�����ɿx�B������NÐ*�q\� �`�F�;!�u `yCuV����d�<�o\&��|ֺ�۱O���"�-�n64H �i�k%�Mu��?�p�<�i�]=��eN
 �O2�6��M��.u���\o�6��W 7)~b�4'�� 1L�T�D�q½|	g����k[�;�5P��woOԄJCTUa� 95l/�pOOO�WML�x�jj���'�@Y	

�N���Lx��+��|�~ivu~d�r�ӣ�8]Kztt$����ʂ�<S�|�⡾�a�d�q��k���Ol��n� ��鰀�m�Jy�3��NQ{���:wySHH�<��S�:�׎�'��~����G@i�@p�ڠ��2��+p����`��' @���s�t��x���∐�?��
|�Dg�!!!!?.��kiiI�{���������###vvv{J�x��XI�I���Cy�]L�3��:�!�����{��w�^R���t�sHu�1@��n��c���6�o,�� �"�ʝ.ƺ-��7?a`ce� �y�;������L�I��E�7#���o�"�O{:;쟛#��.h ̅S��M>�Ԥ��]���]���O�:�(������ 
yU݊&y�r��H��ڌJ� ���c�7�^��\����n̿�n�y��s��]ZT�;Q��� ���ǘ��M���������B�N��2<f47���d�]>�]�b�|���3���"�MTK�X�ȫI�ɀb:��=��0o����P�i*�b8LJ��v���5+׃�Q�a�󫽩##�yHcmw2��� �e�U9ͽ{9��_�x��Ƅ��w��Srlw
S+("N.��O�d���5�7��gƋ�R��O����f�L�B����"�_?g1^�G��/O����z�}_�u�����FKK+��
��UUE���ӿ�	�e|���Բ]���/$�y��}1��5~�/ss;v�oÔ?� �V�5��	��(��F0�Ƴ�-���N�J9���1~�M �j׳ck�ʃ� �_9�|�k�0|�ޮ_È}�Z^����C�*kш=`8G����ݒ��"�����]V��@��,&".�Z�����PU=_����DD��P��.��R�S�[�������������Z�z/�̙���93{���\�(Q���Rz�c���0a77�����x�㎺48Ȁ$��T���IS�����o>Ck5O�vm��)-��(����g��.)eff��#���c���������2_����<��968� L�(�^�y���a*�k/��U���p��p��qqp^`!�������k\���;�z��84�ZT�C񇫐����f����%@	�\[ߴ��M�zz�f������+�����0<��d��Э���|�"*}�m���aRE1d�w�����nxr�k_�>��d�W���A䅯����傞������zK�|�dA�(�dA��oco{��!JZ� d��A&���%���e_�g ��jj�jj�NvP�����T��j��������/Z�:��ڔ�����'�ŅtXeMP`M�������AiU
�T
�Lv����oӲF��j�Ѭę���85���D��22`BWm����$��R�c�^KA[h�ϡ|��U~�]^����P���JR�t���8f�غj�)���X�ҩnW��3|�M��y����7��HfSQ�����o�z6l�44֠���6=��c;�I-P�U'�j2������|#�:wu��j_����f���@�W�x��΅����41;�A�s5� S�x��H�"+'��?r�R��z���u���<�?����=�A�|��gG@�e�&����N�Ƈh���?{��k?'�����v|U
Cϕ�+�"�����58�c�X��Fp�|A��:�a2D��ԏ��G��B��#�WNOO�%�����|�|KB�/���ȣa\�����[Zh�Y5�I�5���a��2c�E��e���rV����3�ű��|��bvb�h��&�����Z����	�'���ֿ�"�IwW�Ъ� @���	>|�| ��Y���\�a��c�'gҹ*.���֖bT�,ϩ��0��̀8X�S�o�����j�:=��?�iJc��#��X/�-��,�װ��[{s=�̈́z�
���������M�$�%�S�1Q�7���Ǐ��K
�>r��2���"�32e�������֌+p�������7�2	�y]����KuJ�J>T"@�(�>䨘��F$�����
O�W_u=�-���q^�A����"gg��ow��l�&RI�+TX�7��K�A������}& ����"�ST������%��b9S���������G�{~^Z�9>p�B�Q��	 ����D��9??�S�a��"�{�4����̈́�,�b��}GH8`�t�
����)7讛KLL<��W2JW����"%��$�vz���GW6U�m�������(��~�e:	99ƿ��-h?1y� %�&�� �R����'��2�Scȍ�팁�b!e	�4
B642ZYz�_����i
��%�~�7SyuQ��7���`�~���%�=�F������}�&���*`�9�|����|#� ��M�&��>)F��r��m;$p)̀���2��;8���p����R6&T��ZĦ�y�q�%�(�Ȉ��D��\�"E!�� �(iyy	��������Rε�V�d�72�����Ы�)&���Ã&f ���o�>��y;L��"]}KK4�z~�ۑ0I�_�̎��~ �$7�F�T��X5����ԃ��t�ྫ������+Zy��ď@�����U��5E���̐�[kJ�}��rn��	����R�h��%��{�U/]�.j���\�16].��w�S��;���X7�1U��.9-yp��� S�L�ͅ�6��-()�TP� l�Y��uȯ_,P���~C��7S��''�%-�
��^�n�[��T"
VPT�}i,����Y��sT������T ?�DyErB�-�ZȘ�P�.:�/_�u/E��� ������S�\���(%��s�o�ao��Bg�h��@�'��������9�/�6>���]I���<���s�إ���0y5�u�L�[��O�1r����lܫ����*s \�
#�n6��e�y�Ԫ�
� �,M����9>�˳mh�S�+[Q�2�E,+Z�&�SӞ���<��rss)S3��]��o��.m�\ _�W!-#�x*�+Ha��I�H��}`��	8�<K��	[�y�qe's6�Kt0Ґw�L�����LOlf&%�q��d�m�EHD��x��%%�?FIM�����������]��k:���>��"Q>�߀�by}�`h����UuT�M��DB�6��S2��V�np�\TTT�?����>�#k���y�����k}��X�w��!+_����i{S�/�����U�(`��Q� �h��(���b3��̀s�~�l骋�85��hp{�����?U�ix�\�����B�%1 �М�	1�9qȶ� V��k�� ��mlء]Q�����E퍀K{��/M��q������}A��﩮��C����A�Z%T����Z0"]ӰAC��aqn��ֺ�Ճ���#�2��S�r����i�;2�xM��H�v���[�TD ��������;-�
�T��L늃<`H;�.el��4l>u.P��!$�ҶC_t�"�����@�(���y�©q�!��W����=�N%C�������@�wcB0�ɉ�"�����MR[� ~�� ��O���;8��|��I��"����QK+sl��3�w�چh1U���$�7�!�gw�^ɵ:[�d"��{����p�F��x����0i�!�a�s��������n"��.�.]��.G%���q�����]�o'��ˇ�]���G�B۠�$=;&=����yX
\�!�U?̓���������Ѣ�oz����J,#�!Ĩ?4d������[5��d~��g����}�m��W�����7���C̊����NW�S�{����Ǝ֎����6UC"�kh�g~"�#��	�E.��͈�b�jу�1�MA׏���M�h��%�$]##���!�q�Q���;^�h�Y��Y��3�$M�#�A�"�)��j;�����^�_�vQ�|�~�p}-Qpy��}���K��]��T؝���ٴ�rneF^"�A��|ù����?��eWc�;��u�2����y��YYY��qy�=�0��[_7\__�Ui[\$?888:=���<�ݦ�
X�l�_��M�]��7[��7���0S�q��Q�x�{vF/����"2���k-##��G�
���q�a��P�X������xy�jL�������`�Y��;���aM�����w}"�A������r�{��+t
)�U���ھ�#t�,̙&��^���T/�HdU�Q:*���@��@���'��4Ʋ��Ӻ�#��f��/��n.��/�C&�+���¾}��������Q�-d�l�>�7��'�����	T���Ʒ�F��B�HB�p[���p�Ğ��Y��|x0V��%���G�V�Pj-aL��'��K� (�� �Z[Y]�lN�|v4YV�f(G��GQ4��1AR���V��\�h����6~If�wd��o�ޔt;�,FL�����.Վ���=��]��|��3�#�3c��z�%_��H������~����W�	8�~������f,X]���˒�G��WUS=Of[�	``U�klH������M��>ⶼ;�I�5�p,�M��|�-�}�@�^ʓ_;���n(RR�g#��a�O106��g��=�yd d]i2�cዶv��["0��R��B�O+*��7-�����^���#Q&�pUK��!s�l�a��	�Gy��M�×�����Y�?4���m�N{���I��@c>0p��ѓ�DErw�ȈNM��A��_.�o�~HIҮ��:��iVY�ת���g/ B�M7h~0	�q�M=�� ���	j��S6/�1v50�v�Na�ЦٿH'��e�8L���*�F�;v�Fhzw{9V]&����O��׽i�E��Gq�'��]+���K1���^":���婼�X�/��th�����J���aO2X�M[y7M�w�A����Hnw{i$��T��.v�[A��4�z��F�ƾ���x00��qu������GO��AV1��G)墉:���������pED6�Խ���ͅ�#��� �h�n~���"��ӡ���P�R�J����9��C03-�3,Sᄬ�Ń��@���%�)if��a�Mx��i���g��$Kf��9��PPYM19l��^�'r�7����E��g�_�!D�;k�U�R%��6z4��6��po�]�=L�aK��f��s��lwO$��Mƀ_�"��+�w��=v�5�n$��m&� �����F�����Q�������XP��]V��q֊��l��%��l�Bv �ڼ�Q�����U^������9zHQ�ϊԘ��
�ZZZ��˳I{gY��^v����3(�h�@�s��Ku/20����#�9�<uVh��a˭�[7o�sm���$`�bz�2MSǙ8>o��M91ߥ���uo�$h1���,��_���& H���ȥ���^YS&��rx{Vn`qc0$?��&�@�GY��w�c�u�r��^A��U��
[��F��t�e���^=c��R=����'�����x1��Kpq�Ia�[�iԾ�\F��sN;�l�G�d���V�u|�ɵ�4�tJ'�[Ģ�WT���m5���8�u�4C9^��E�Q����gj\v�*H�]�*-�� ��wFJd�㯔�>�f���9�u�I��3:�g���Ζ������ci~k%������b�T_�8�������K&��#I��&�,��{{�뛛?f�)��o9r��B>��<U��EE��xZ����dh����^�ٿ�Dw�xd�qrrr�&5M��MTĵ8���裀��D�9rwG5߄�]��3�_ul>N6W���_���Pݐ�v�=S��R�'�G�3e�Fi�������*�!Q��ki�h^�������~�Z[���c��(�K�p�C6���sb�%�E٬,ܨti���ʷ5���F�r�+����.&v1�7�mޡ|K�����"q�oo�U7lZtX��� �%En����1�t}C��k~~>53��6gw�G��y�ݪcʢ3v��O�zQ���&���x�x�
�.����B��;�����c��V�ӯTx��W��6.R��Jά��Ɣ]�ؾHu��'���W	�s�'cg,$R�NZ�3,�h0��s�-����w��/�+�J�q��p�'�y���z��%�0Z`���Z�,3ā昴7�������Oe�Tt7o��G��V�q�J���2���7���ee���ճ.7�_����� gs�E����7�?��#B���q��-��	vJ�z�ԭ�F��҃�������=B�2Fon�?5ge���HL4xU�F"�a�{�LO�؂���3�<#��C�W%,�K��G��.o�����f��+�fJ��2Sk���πw���x��'�t?���ON�)l�xR-�����~�nל��C���~�Oc���k������N�SsM��pI֋6�M��Vw+�X�G�|j�wvȒ�y���T��K���z��K�?90����_����lI����ʥ:&ߏQF��T�[�7ܡ�D�>�g�^�&&&4t��O1��}G�������>�te�X�臐�����|"�d�����%�w�İ�@o�L7q�/�S%����ْaY<�O�}������~���"��7�z����TD�	���j��H�hS,����ˮS���3��8��Vb�o�H����X��5�P�O��<��z���m���h���r�����}���t�q�$]�K�&mU�������8��fgF�B.��k\W�-�=>����al[���g��L�Ǉ�~������d^tБ�[����}3��Z�+��M׼�>����-����Gi��[�S�m�x�^H��>�4��|�{��S�\ht3:))8��������a� �[���Q%m�P��V.���H�ׅ���OR��bݒ��1t�Fo�<&z�;ߝ2:��<n+�����u.���Na��M����}�!�n���ۻZ\\,�,�
��K��ϯ�)
�B�W�&�����`�77w�ϴ�=��6GggoH��lk�o�*͘w�5Q���j�ˆ�����co}g��ϣ��c�Y���mB�ˠLb�p#��j���ձ�\����������Zggg�_�q�LW�={��o�}S��������5�����T��ɓ'��Ъ��9E7���(���FEGkt:��t�U�:�/JJJB�/����ޮ��̈�KHH��1k|]���^����'9W�O�/6�1j'����T�*�Q�U;��IƋ���?�g��B��㣖��B����h����X~`h�%�ǰ��7���[�w�2������!r:���$<Xj-��QZ����K����=���Bc�H��n��Z�P�|�[��F�5�_���zܰ��Lƥ�޿k�����**8����w�k��ag�s�|N�_����^��������~j�M��AF� }Ť�5Z��Ns���Н�ҋ�����y���XF[999A�oq<A�w��y:�wwo�����^;h*���6++��d�|��#�wȆ��r��|�i��t@����c� �7���w�ߊ4J��qC�n�梊��*�+�����v�`}KH �z~���e��kE��y�����C���%EΒ�����)���^$M~k5���sO$���췐T׋� ������m6��3bA�?��&z8y�_~���FRh���	����!�iq��6�r���P%���h;7���f�;���;���~q}}J`_�HHBzz�S=>�<�ӽx���ٝ,������������n�C�7�w���㵑&���k�;������P���r���Iϩ��B����ӭ�嶧�S��Ħ+��-@��%kW8Y�g���W�,g;c� ��m����DS���J����涶�3^���jT�̨N����Ϡ��{��HI�&��3A!!#���*���O��d�����@�@�K����!%~kYP�V��7������ݦ��?��(�[W'gg;�P�Qh�K��"6�Oj��'rh��X...Tn��'��Ç�SG�w(k;;A�v[���3��О�Ga���o��7αY	�(����W���ݠ�_�������+��t���-��!�uG��{���՟&@�!l�gb �p4���We�:P���\}��pw�nhl���_g��Q�]����k��Lڳ��O�m$�M>�?͞9~��Z���R�F���K��	5m�[nY��
���71A�����'�^� �ǰ_n��y��l���]�!N4~�?~�_��R���]��v'ԋ����a���б1��$ev[
�WІ�@�1�ab`Ў� 

�������T=Mo/���Γ�Z.��Y4�C�wFs՚�j�(o!�fp�����s�~XT�'|s�o�v#NJyqqA�����'W���7r �K�Ϗ���
��-��#�-��)�0^
ll}5r��{�m	�r��>�y� �L�xޘ��Z�`�T��T2���a�DH(�5��z��<���Fs�rR��	�Lֺ�|׸g���܈�X)}�%$�=n���8�H��x�W*tw�}� �D�-�uf5��|5&=��T�ǻ��Z�n���%i��5d|�j���� %r�<n���xxy��V�o�ٵ ԕ�y"�F#�1?����C�B��;"���x���̇����̗Z<$g�XXh�#��/��Y�n�c��|�H��B�n���u��9fcy��6��R�Ku�^78*�~��,�U��2?E��"%Sÿ���z���a�l����;a�#R;��&�H<�"(�� �e�ڑһJ�ɲa&6a @�JdH��d`�������3��ۛ������<����S�}̓O�y ����<<��xLr�����jھ�@l����0.��T��!�:"�5 L�|���]x��W^^����U%�pe�]J��Ze:"zB������02>G�}eO9i�W��J���z��tk��g�1�t2�66��"ȣ xI���W'�|�4�<��W5!n����GO�kfx||���J��ut��29�r)��xew�&�A��/���ƏY�����NW[�3<�"ۧ�g�!��I7��!	��Ƭ�	�>�(��QdV�ٔ 4"���!#"������M���o,?����i-�a���!��~�[D��=]��!����t��@S��ii���1[��� (���PL|G��&���Gy'^=��d��=�{�Oͮq@T�Z����~�!#���0:6&aF.�:��؋�3X	4��Vհ��p�î��{[ �o[	H�ss��^gj)�*U���Qv�S�G�H�e4x�O���7�2@?��	�V�V}�;@�k�@��= �d��2��7f���R��7����;���DFb�|
���OቩXY_BD�OFZ�E<�'�jj�w	A�������x���d����h<ł����O�|�n��$Ϫܞ�%jܟ@� FFI�P��1��沲Hqq�H��ع*����6~���`��E�^^�i����a|�}qP��!�X���ó~�ѷ"���M�� dT�U����*|��B�ו'222؝���������P���F`
O��Qakph�d���.�ᖟyK�4?��;��~v��^WW����']QYY(k�k�)�N�R{ *�ONpf����=�*�2��!�%���tT�P@�M�^�q_I���zG�Q4a8��Zi]s���lc"�+��3�&�G�1�*|�1SaD��Ml(1g0�N�f666�9�I�RF��W���t�T4��f$��QL�tt�K�"���~�E@#���{!w��FQ@z�}���Є�K/mj�@�֒0Q��-��^������x�& ���ʆ�e���hh4666Yo�]u|�PR��<��\K��������uɾo3T$MܳЩHW�btLL�i �L��ϓ^�$^��ùZ6���N? ���D�H�����)r�
��Ĺh]5��bGG��������6 �輝x�oX/���I��O��ދ��¦�	�խ-��G�mFF�$`�^�4�p@5��zc�C,�P� tD�ꕿ�}7���c,O��'��gѮ���������9��F�vy@{�9@�%=#��۸ۺ�������Iv�4e]B�V�W�>��<��@Nj��prqi؎[-48��	�?E@{��z��j#n�dql�̻w9�c�) ��5�����K���_1@2 �>���"#!ed�[���g�<��u<T�A�h��H=<x��L����c��U8��z/��ʊ,H խ�4�����+ռw����Jv�߿g�JNJ�i�<37'7�Wk�������Ll�Y ����w�U@��6:�'dK\�𻨌�@5�
*b��h�D@�_.�gff^�MoF4+<�r�u�L�4��Dv�B`7�Z[[~�Ɗw��`��@ᙁ�����"#k%#S�$22::�X -�*DLr<�����c��*|����C��̡s��|�=wWL|����|����t��S	t�W��3����0)���w9�5C�9��ob"L���3a�u�KIKŌ�'uhzD�Sp��*ъ�^%&��0��iu��L��ٍL��A
A��҅�~k0d����g=ی݀�rV@�g�d�u6�u�� &y՟��P��^H_��U�)�1f����RN Ê�'*���v�k�V���=S��듍�X�La]Ȼ���F����i'�LAQmt�RY�U�'�d��cq���W�U[R�J�ÓX��(7�]�%�n��bg�j������5�-�[@,P�Iqw�Jc1
Y��G�!��ss1@-����kJ~cݶ{�� L���� s�iWʔ�OE�Ĥ��'�N=S^�C�	�Jԇ���E5[]Y
b���E5n+֔h�n:<��|E��W�ߤ����y�=-8�y�P��r��Tx
.k�dEԧŨ�y�8��ȵT����X5�_e1��v���K�)18���}}!�<��(�*����|���I��dde�������Us�{�Pseok���?�~�G��VO���̧�1*+*�Sy�mJu[:'�}���
>d�+�p�,���m��'1���������'�AbPM[�~���N$��������2�|�J�4��v@ܼ�����b�ۖK-�Yd�cc1W��r]�Qa�{31(�x�s��3fs5�b�����U��"W:TmTUT�J��,�
՘F,ٙ��`�iD=n��?���(��K�y�H��SV5U���0-8��UԾ���呔I�|�N�N�)sP��a-�_1i^�jjhh�<Ҭ,U/�@��\h������&��8�S�Q��r.�҅"��t+��J�<���X�@����d=�;	(���#�H�W +$PC��8� K��XT`��k
#~��O�@���p���y�tީ�N��<�t�ݙJz��̙��0��o:���i99�?������)�S�fBz:�z��f7'��6D��SD���%O�J����[@
�+�L��-����~@>Y�wvv�O���U~���C��P��x�Z�d��E�Fix` R�ŬE��@J،��9�$ H�8ދ3��M���/Ml�i�+gK&pY��<�X ���Gcw���z��RKH�p(&�K�L�����>gkjj*6)�E9��E�
�,,��ZwF�>nW���o���=O����k�}��611��מ��� �$��\������}r��?�\���v���Q��ŵ�?�&����a��&�!�i��?K-3��@����p8���g��>�8-y m��9m��Ag���R�)���u������;��#�*�	YiiaO�C�>z� �������6�_a<F���8D*4 #����짹U����@�-J��y[Ɔ�>"������B���#��]����6|ōG[Y�W�>��%ҙ3L艩<��H�]A�h���SS�e;�F�P���:zg���+�w�FG�1BJ_��hڬ	6���μҷ�(��A��p{; ��2%/|`D&�'��� `�h`P��%��Og�3�n�����O<ov�4t=h��Vd���f�#��,HG����xnL�������Z�P�h�\����,�>ޗJh�X���Ӹ�6��=EP�mPG�����aR`�~�Q�,1wxG_<�h3�ׯ_���r�뉢��� Zg�m�45�q����x�[���(�|�2:�����w��q?�)����#�JT��d�=�����;bl "OPHH��B���D-���D>>�0ɒ N� x�W֋�3*X'����5J����� �,��W!�5�T8i�lr�p^�0�cv�C�8��љz��ɒN��٭�~��/��[A���g�1I�nwm�ڬu趶?S�r���F����-�̓�?=mm_o\��q��]�:^��A��t�WQ'j3��[M$����w���|��:�񳜁HΝw�������P�G+��/��|�KE�����^{���cV�M<O�<ys�|`h�ޖ���8<�.�f���n�����p� ��4Qt�p~���SH5-1����	�F�������� G).��#�����F�|T��<OxH��k��7���/)�+Z�Z�Ko!��qiʃ;@KC5Š�c Z���>~$v�<��
�jv���c�V~��[{w�T%TU\��ZWX�ݖ��Ŝ���)P	<�ׁ	���h���U{�j>�:c=��ҡ 4ΜYe`(�kG�ʾ_�V+�8a�f^��o�BF����4��D'��,�B�lx �9��{������,&E	xu��GzLHjALt�/ �.�K�n����R�.�2���[WG���:�P�oHQQQ���1��̟���	h�,��|_��}b^Ml�5����CȤ�tt�;^��,�D=9!�P�CT�$n*L�lj���6@՜�k X�00X�#���j��xV2O���A�tq{��ـn��Mi����q��V?���b����_�!/�����wIo���h\���|�n�*޻�⬛�K��Ͳ�|�=�}u��.�'K������5�H�������Iks֭{�����I�j���-6'?�:�z,sȠD���
������GΌ��tF�LO�DH���/�z�%???,���b���dU��3=Ao.$��5�oX8"H;pzOd�Z�:Ma�g�0TdJkl��}��E�(��>Ǌt�J��S	ź<�*�Ű�����?'==����(BwGO�z׳�VL%xK��܌ML�T,8�-*?��`_��<�bⷍ�#k��Jl��,���<˧<��p	����.,�tv*�����Ơ���zk�.m9[%s�����Z�,��h�d..��3�׸���y
�=op:L� �����/�����t��^��+�=,ljj�zu�_e6&ig���%T7ZƱ���Y�"��߶P��6��!�B�x��29����s���rB��-&����n��n���ׇ�~�8Nx��֪PR�v&�啔�j���T'�~��mf�#x�%�#@�{s��?����
		�p�|c"Y�$�?ט9ɉ���[��c
����͙�3xx"�FIٌ�xx�)������r�B+���<#q^�*���?������#�bhci�`~{�h(1��e� a�m �
�.Zn�1���%}g�M�`�ndl�2,f�]�$���߇=Uq2�'u�jJC�rC̊g��D�����&���`�X�Nu�b����ȔU`ӵ;�n �	���ȓO���l���ڋ�=Y�̰P�x{�z����&;gWW�q���Í���\τ���Fi� �$Ň����'����	X(>�����j�@�ajYS�ov{q����\��֓���3DD�����f
�P��@����7ѥ477�U���J�c� �癹C� �d-�T�k<,�ϗ٬I~% `�Yz���@�ȱy��nҷV�4����y Fs�� Z��Ѧ��PȳIB*�'�P�|��:bL2"���$���~��(��˨�Go�.��C`��bgk�Bh�~�{��z� �C�^�1���OX���m����r�]u���8f��<y���k��嶤�Z@�)|N%jFH���SXdda�Ԓ/����;;%8��]��z�|a��*h���)]�0�̈́�m��ى�
�������F�bCR����|�в;� SS`[�Syu 8���F�G#��_xNY�����<E\]�I�z#$D�.Z=o���@�ŝ��ǪaR�
Cdh���[���B�[+b��sw����Ā����qh6{��
D�oh�: 9Uk@���[�~J�c[X��F��;+��R�+4a���?���ð>ב�D{��d�?:���f0%���1T?n 3�.�KU�dD�n2D�/on��� 9֜�FDD}����@D-����_��X�.%h��Z!���������G�f/?�{��'�]z���������Mqqߙ�mbu�������!ϳ
ǹ"/..�@�r>���6��;V���!��8�C+h�ȯ�Ȩ(�3�O��@\+t_^N�0[����Sj���ߝ#;9=����Y_@-��]�Q���:��t]�5��EĪ�j<�d�q>����]�L�8��+���2 �Ē��@ �2�:jj�ȸt�`0b�:����@h�/��e��(�r�C�	ڨi2#��B?��sU���Rx��O�W�;���i�Y��/�\`��=H_�9�R�wA�G
��Yt���a$\e��I�r4o���k�!N}��A��2e���@��z�&!a����\�M��F���*�#.N,�_����>��,=�����p��[=8��,p\T�>NjY�4_.�v�n���daH�?�MY� �=]N�(:Z߯��� Y���h� �bw8����[	��W���4����xW:�с7���H��!������w�+�a�����Bp�z@J�.4pN`c2�,�r�Z(}��V~xc�P{���ݦ�������t��N.�[�����<�6��7s�����
�8H;��|R�._�H��_���tr?X2�s��c���Z�4��W��,����z�H\��fʰQd�Io��ZN�/����_&�p��WQQ��QG|�T�g��pm[N[M�f<00 ��u>SiBuI����K�x�OT������Bm*b�̦���4�:44K�ru�]so"�~���i� d~7� 8�Qh�).��bJ�,�T�^�D��q_����o�C��{)��&���q�?Ť�)���i@%����X+533���.�˪�U��p��&	S
� ���xS�P(sYN����Tn*B���p���� q1�����|UT�мA��33� ��Q.�7�D���46ŝ� �4���5@��"B�� �	 �ށ�	�ޡ!z�<C��pgݮOr{�_�Z-4ġ4ZL��ʓ��� ���ֺ�4���0����1i��(<����q��Y�A���%��9r�js��/�hY�^������db Q���eC:Sa��_��!���ƭ,�OB"����
::���KR�zh�a���g+&��?��7N�W��zq|'zxZ~���o,cn����^9�'�j8S�]ߦ�s,��p��'[��4�y��9��On��AS�iKu6��3!�l���9NGI)�o�o����B�1V�����Z���f;%�m�G���D�T�j t��MZrrјP����Ύ$�E�����|���Nn�n8Ϗ�)���c�A(���<C>��c�Z�qĥ�p8�ݕ+Ѯ�������z�#[1���'J!�7J, #�bWn-�m�i�:�B��?�2ۧ��bP	X�V 5�`r����veA�pR�7+�����y_�P���آ��=LP=hM����0	��%����,���w;�ۃ����cK QB럌�ίw`
ź#�T+��8��;���q{}�kԟ?�L�ll�]N��g9%2�\�Q�-�"x���J3�\]�����\���j&��?���g�j���b�wGP�J{<Y�
�ٛ���#=���o� �Y{Nnn����Ϸ���i���y���Q��%�Ĥ��s��@~񥃔��0��8���<�l`��5n^���?�泘-���2^��>��ɺL�)�.C��Pz)�	0  �R�g��uӅ�h��p�"�pjVVVr�'~JƥG�2U�%�/�>qsq��"d���5���kkk��נ��z�UfԮ^'ɭ��=��������ӣ�~����V0^X`��@�gr��S�\=$�h˶���5�͜֋)@�v�I^�j��k�#�א �����?6	0Gb���K=q 0��C�9~��/���W�O��k������ .<�	�V1�yn�7�^�~m[a���vkdU��P�'mm"g���i�+++�D33$窔�&�����𶁹�TR�,�����ws(]w�/9�t'��v|N9�O�G���+�'�^���B��4�@q�$q�1ى����+��+3���k͟��C�B  ����4\�iD���j��+
Ί���`*|&���66�`���}�������	q���Vn��/<2i�%�u�tAYNc�uAۇx��7���ߔ�>��m�b�����F�ɐ���h��e>r����j���JW[��ȥ��Q�P���(���Q�l�E/�^�K䠵1iB^
��aL�w�|�|*T��F��L��)�)�g��\�~x�;�����+%\k�jӻS�1 ���b��<�s��U�n�w�r���K��#S�۾�'��m���XlO�sQQ}��.�X����m���ld{=>��3�����\�f+1��p�*�����
����<���JGGg�|��#��aw��&�uЉ��S���onn��Q҇�o�EQQ��lG��]�͚�%�����N�Zt��Co,��gJ0�^��;�m�ʖ��+���1�@s~�XX�^����C�ԙ��Y���R�'/�%$$���XDR�Rȧ��; A���`��.�}�kC����ӡ�W��4{{/|#��S���iҁ ]����p��ϰ?���l{�pg47뭪��Ϻ%Q�6�/}[��-�C�5����R��z��p�,��ݧ�-�/��f�/�P�_ e�k�����\�z���Xw�4 ��<�ԟ��Y���xa�{�d���5����+���{L���4đ��������q��4~&�iG1�M��kz���B5�����J6_jj���Dl{1轘�O�^�ے��; щ�bO��&逷��ƼAd���ϸ�.�g�$��_�J�grn;#w��X��^����Aʗ)����QV�����hn���+�u��B�����	��I+�Q��Fd�A@��3��7�S%�t:@$��Y�	0����s^o&[�O��3V�$ W�����eD�3g�&08���;z�����֖���~"�$D�Aƭ�NWH�䅃�|�ԕ��dal����?��+����Ȱ^lJD���� ԰�w|���7���(�@����t��K\�s���:"(>>�g�b��l��,	ԘՇ-�����`T����ҟ�6��������x3W�7�#-�C7���Cyi/���+����M)�#�C�������$_��*(`T7������ja��Wl*X��}�"�Њn��h���W��Ł�f������J���۟�d�VA�nO�R����H�s��c������~�����u�3-�'حvp�+�Thli���`�E��ҧ�hs'v���y�kEnrrrP�Жl��2���;�}ꌬ�]�RG����44Ϟ"��r�߬X���;�k���Sw(���2��\	���C���O
��]�Ɋ�ͪ8hVw�

�_��i�t��J'�aD���@�&W8�e�����^�].yIm�_�Y˕��bc�@���� �d�V��������`x��_��S��k�k�H��m}���LL��f�zy��Xߝ���]�{��s_��?�ۮ�N�*�(("���DBA���-17��z��`9��4Yy{@���tt��B��H Kv�|_���W,�L�ٕ|�m'qp*C5_����ŌMF�9�2�=�in�D��Ƃ�t�`�򑋋���f$PW�~����x���xaL��O�5��F'L�����EH��5������Myh
Ϛ�{ �#?oD�e� P>o���ȻǼ�C��!�鵇��{�����;����{��B��eK�k���A�޲g��*�-eoٮkvmQB\.�k�Ȋk������T����y�s�u��9�y���>翯5��]GE�j�Ꙭ�T���M�B���Gl� '�G'
~Z_�/
"ᖇݵ�60z4{�!0�)��sס{ ��8������.����9(x/���a����� �|38x�/��Cu��������YE�BW�EB�D�v�@@R2՞xQ�W�����,!��*�:000]�k�*aOq�]�=���
��TY�`��-LKc���*7aiShp01p��1����8���@�"��b�����==�%
������A::qެ���9�U늇�	W�	�Q��]ZT�����F��0Z6k�--v'��4=3z�{J����q�Ak]���k!�ׁ� "!��M.I_�x��x����+��6-5`@f��D������cN��OLN^�ї%w]S�AZFF�2�<Xx�A���O���'O�g����������=���C>���~�g[�X�N��A���	�z�Zv�5������_g�q2�B�Ѐ��}oo;�خ�ޒ�0�����^�)�9olx���������	)��N2�������޶�=�"2����}���OCF#�G��T�W¿#A���n�����U�Ԑ����G'^f`q�C]w�X����ۄx��2�Ɨ �p�	p��k�	�\!��cwѢ��W���}�,Jl�%�!�I�IH��ߟ����~��QQq�9��_�$D�����Z|��C��ҨB���)'�i�N݈Rhd�_X(p3�����Բ��J����;w���$j��_��x�˰�<����`iP>F#�穠 e``�+Sr�\�4U�����*7��c�R�aǲSs*lFk���f�]���e��UH��i���o��;����^��h��ŌS���w4�����U ���mAf�����廐d���V��'��o���!7͆O�E<�ǳ���FC���K�>�H~���P#�՟K��������P�MR11��,�TU���g�%{��;'���w\��q�$�#��ϡ�Z�s����A��C�<��!�M�����?��NT�yM'�j�_+�H.�+~���kԕ����5Y�n�A�_��Rr~T6���݆.�����o��\�2C��[}3�J�s��߿Ia�����&��c1W�Wi�<2���`F�S3�N������d�L<޳h(1����俑#X�b-���;����..."? w��BJз`���}u���*�N�b|z����9��� V�>@��43sfqE���i'`3=4�&Su�e�W+[ۧ���j�~�`�Jާd�k����T�sVFf�b���hfm�Y�tJJ
��*{����K���k��.,����.`�	!��J���{̬��e;�$�VT�sנK���q�b����׻�ty۾D��F�E�a�2{�ɻ`B�����O_}�ޮ
V/��Ą��2;(W��������]qTU�'�LE��N���V�%p
��qʾz���^��O	��U-�ͅ�/^6�7:�1��mu����e�P=3���6��[���N��YJ
o#.(��Ǐ\�Pʪq�~~*�9|�*$����~�B�Of�P"����=�H��`7	�߾��	}�]�Z�f��&g�s�����_z�Z399y��)����9�R�V��l�9�[EF�U�R����ssq��|�N��|,�h�e�/�p���z�*�d{;�TQ�joeO�W��$l��P�&�@/���gfƼ{�$x0�ry��/<��04�9:9�ZK=��a���mW�F�J�~�MJ�2��@�FG�)YAAav[������G��gj��4�s���̘�6�|�"���EG�Q�]��8\4��A��/�x࿭�����s�#���Qc�(�QM�'��Z[�����1������,hv�	���K��x�s����w����A�P0�T�0zll��,i�_�	D�˧̋�%Zq�"�����퇧�9	�*�
dKt�c:�Y�{��nnq��W�M\]/�gdXWwEn�m3������>'�.����Fz~z�8�h��#�1Xw��ݚ����g�(����R�"t��	&�/�>���9�����l��b��~8/�s�a�F���`����[��c|�Lt,"
	��bZ���٩�8zB�=G�5��w	9G���4;���M��`n��a"������f�d�:z{i����lI(���Z�qXDB���$��S�*��|d95o���8<�$|�X�Ei0e�	O�ហ�CB������@�Q��P��e�5�M�N�,���Z�[�˕F���(�]y-��&�F&�<5(l�I�BZJ󜂅�d�=��/��������X�E��X�N��P�w�~��J���@?0.��� ��8~TjR�524Lߊ/�T�Nޟ��6��\je8�@޶�;����@�`�h�b!o�1�#l�� �/�w�����NTN�*�]�7���B�������W�9�:�+8w���#�P�Sn@��/�w�0�c5�8�J�J�������W�7�g�W[|��7���t��c~�wUv�ڏ��?�w�؇�8j�o��p����-FA��J�f����b|��/���|\�O���@�? �W��m���e^�_�@�;�b�G���'ֱݦ���0G7u�vTZ�a,U��`�.D3�c;������~�HG�ev�Il�D�l��
����0�w�%p2}�ۭ���2/J����$�nzDfi�F��y�z�<��ۥ$��E�݄���CЀ��˾n��3_�p�Wn�o�����t�/�������gb&J�WS�W��򒘁V��pV� 	f�W���/�0K�P�"SX����MDx )\L���kf�o���S����Y:42�ݼ$q�Zp �[<��z��J�{bQzh����)�X�*�����qӜ���d����Ғ���e�!����9��L'�Q�b��5Q�ȱ/����L2��A���:��?_��?>Lg����S2�������=~���t����� N�����#���.����� yi�N��I��>ۤzGM�5w�,7��II����O�>B�D�K-S�j��*QwF�,��@r���ם[���o�~�!�I^ggg��W- td|�m|�UHH��������G�G�)��g$$��_�}1�L�W��֙�E�A��Z^ �	���ٍ�$�C	0Z(�Ũ���kB�nl�����&J'666��×*�_�>!����-]\b�P�R���E�2���^Cv#�����MN368�xJ�<���"��U��n!Ϙ�OU3��	"\?p��h��E�m"~���j�<T�7Ď�%�����2Ggf��vR��iO��dY���Ѱ��P�uj����}��F�S��=C]1��d[	���3-Q��jC.��yg��=�;x֋����拂��0��^(ҽ)�5�������>qRb����������3WlU�@�.Ňߧ£!a�b+sC��9����Ӊ
�;��k]��I�+S��<���*��K�S.?�r�!�++0g͑���(�}�9�	*H�@��$��&D�E��
գ0{L]S��	�EfP<���-(�@�'C!{あZ"n/�lF3����IW��y��:���}���]��*�x�j&�o�1g��|=��%����n�(��*>�0�OJ��XMZ��U�OyXօ�+ޟǜ}K֌�R���ܸ��,�r����ڿ"?�z����6k����@��Ch=�A��C���^0g�C���?���V':���fF��$#W\]C������8_ђT2�Z�f����W���/�)�K���񩸰��w��^!-���~�rb\��Oʻ����̫�N��;��ك��:��B��K]YhuK?Z�/_��Eگx��-h������.�r���;��
���K��I��\���7s$�D#O�,�yW(1�$�-ż��c�f�p4��ᕿIl�'om;Gd�T!������#�+�	2Z�60Lrp��C���
��s�	�gP'F=Lc^�uXx�gf[V}�
_�I}�,>G�+5�"t�7�F���k�@� ���M�.֏�ȓQ���.�³M9����y�ٺ��ɂ �(��K��3��}<�|e�L�d�1&��/�T"�z��8��@����u�r n���4���'X�`�7T��VP�����GȒH�S W&��m��Q�w��I�A��6os7~����C͐@�:��~
.^GWr�S�%�4�๺�l�Μ�o�d�����5�"B��F�y�~o�C~�jF�9m�6�3sN��^�Z�Dܽ|5�4:1�%(��st�,7�|@Bo�)�R��a)*� !b
1ue�}�h�`�h���#��ʡ	j9HQt��bܦ����;;&I�3�VGP#���nT4�8�+30r�,�!"y,���0���8��85���JTq�Z�������K?j
2��#����N����:���e6:��܋�����ou�l�3;e<��8y-����,�;�Nz;aZ~�g; =Z5q
�M*a/ )�4��2������x8���N��)��\ﮩ@���5�$<�n-������L۸Z4u֤/Z+(����u�b�|�}�|-%�m��V���#!�t�t�im�}���x8e24 �L.u�Id�\+�2���
3�OdA��rZj�M�֢y�~t>0��T	�FQԢ���ٽ��B��n_z(��P��v׉���y�b��3H�T3QG�Nvp�w{�Y���Py��͙�b�����0��m>����epҠH�˵��GrЎF��Æ��TfٰA�!/#����5-q�lQ����K,��R(O��G��|�V���[VFe��Mh���,c3����"Ϲ3��j�O��)bW�e����.�j��!C&<���f}G;����}�@���F�ԱL��@{����e���Zv�1]4�=ތõ�6;2lY����FY����;k���[j��A�A.��6n,hO
k�X��[I��+ق��6�[�5-<=0��C|H�7���ҹ0��&0Թ����H��������쯺���G�K�,<=?�oB�(�M�s�[�q�S���8^�L6z��>]%&;H39�ٺ&�͗��á.{!=%{߿CmV�
�ю�_B�G�L���{���������,]]�ǾM�e:��ƣ����̭Q�5���k�>>#cߞ�#-*UM�&#���[T�rppH���=s{��F
�A]�K�K�Z�!CO���<����w�ik���H���3�m���k�nʋW#�����aoO�K�K��V9��L���YS�c$vA_�}��H׎�S��F�����?:zc�� S���E��k��_l̏��.d��J*u��r���N�����M��ݓy�����x���V�_Ȟ��?���5��[=���5Ԭ��,¿L���>y�e�!�����R�/�M��v�����<�����-��͛�Wi׾�άsŲ���[�
�-�~R�2(�3�8.{?�}���o�_�-����=ſz�1���n���"k�J���`h�����6�Ot�q���a�>�@+I=^���Y}��1�L+��������J�w.�IZ
7=Q�+�kh�hl֭)l��@1�FGGW��X8�f�U2Oe���4)-/�����е�'
0t�/����yR
���h8�SY2=#%���BSWO����C��J�����x�&f攌��I��f>'�MuOO����v�n�Ӽ{���� S�fqH����/z0��6m&	5@q[�����Ɓ�SQQ���=l>�TU�vuU %�eQ�2���q?Iؔ�-@-����.��326����X��;II���#ͱS��y�=�P����hchj�8Q�a�7SO�wہ}G5�i��ΘB�).~g[.ֲw(��MT�::�mmmY]f!������G薻�j�����a�K���,~����w���X���Q3|"�r
���->9�u�Ew	0z<L�F���hUq������h�^Z�T_��#��鎬
g�\W�d��kq�;f"��h8�2� ������
���G��{�s���)���G=ۇ�Ѫ��e^g�V�"����MC�6\tN�l��+>Y��r�~,|�����Բn����S�m�S�<ڣ���3|�]�'˼��O�G��@#����)o㤾E��\�H<��Ul����B�.���8���@�����\�ZڦR�A�MKN~� �Q,Q�٤F��~x�~r9ڋ�����ى����s{��+d04Y��&鬯���0����e�5�v������{;G���M����y���B�];�w�f�V�\��$%�c�@��_g`�qtq�拾�*��H=�Uڻ�闣g'\e�F%����
�0���s�a�k�;£����'+qS=��������St�������Ɠs��Ϩ�����^4;iC��ڌ��հ͐̼� �&�lsB�b�Y�Z��Q��:`(�1������f��i�m����h�΂�/R����)�tV��{�@S�e����j?��>��ǙG�٨ �o�\E�DB��-�������`���# T��B�e����lΐ$dl��r3�XS���y�0ws�������2N-_�\� (�Ru���H�~��|�y���ɼh����R�:Ph&aZ�����b�Jۺ��H`T�y����.WA��3 m8�����Y�L\]��~Q-���ⓛqS��_���C]0d �(�5;�gb��6��	[���F��5�J�f���$O�<Y�A9q�#y��1TqS�`���I@ R��fXT��xGn4�q_��L�m�6x'\㠻����0�ge�$�CU]�C���Q��{����=v�.o\�9&�@�}�?��5�ߩo�>IV��,gt���#�L���Kg5W�ӻ9�0.+�
�z؟ܞ� �2�q�T��}�l� P&
fv�� 8ݡ-
��Gu]��d<+}	݊h�C�)h�{�$h�@�(`4M�{D��r[Z�l3}�=zE�/K]Wx�+�����������cb�2	j�j��P��1l�{ͱ����'(J~�I�ԔsppB��Gr�+E�X�����
~yT�Ogf�׷߾U��z+����ܾ������;�^t�0,�vp�(v����Z�0�x<	�"�v�tWε�0���9������7+���b^@żT���ɻ6�Ȭ�>�ey���>B��žmz>L��Q�/�b����c<���
,��i�.�$�66.������p"���Z|ʕz��0���

��g��.�V�:ۄ���<��j���w[�w?���;3s���/��]���d7���՘�Enk�{��e*��B�E�ylum?�iGk+�3����v���{=[�w?L<^S]]]o���Au]�}\�ԧ��p|QB�������^���{EB���y�C�W�XJsx8���Ji�1���T��R?WGG����~59>�?q�p�a�f4��ȥ1ћ��el���+sss�bcYu$3l�x7��f��m�������;.�.���H����R�NG�6Fj�$�������[x�m�>��H�|�p���t+W�K�	j��CP���nWE�-�|�. ^�����N�3צ�or�=��LӜ��Y��+E�z^�V��z��6tgw!�W������J� �4�9at�>ށfP�(F䤅�	�WY�H��}n9L��LCO/��5��(}�%C:��g��8������1�*g��M���<$s�-Q!,7�o+�)�=�PK   �eX�����"  �"  /   images/a890ee50-b65f-4e8d-9ddc-5b796e5840d1.png�"݉PNG

   IHDR   d   7   ���   	pHYs  P�  P���Dm   tEXtSoftware www.inkscape.org��<  "pIDATx���y��U��w�{kJ���2UBI !�DA"�Jd��->�x*v�zK]�G���(�����2=��L �		�TU�JU���y�o��w�͗�M���֩���θ��9_L��+5�W��5G4�(����e֬Y���&���RZZj�g̘a����e���2g��:u�����Hy�AY�`�L�8�ʎ;&��s�9GƎ+�x\>l�K�,���+������r��Jn^�h����K�.���l-���2�����;O23�dpp�����om��ӵlP���csg�h4j�w�ޭm2m.�HTzz��^nn�,\�P�G�����7N�ϟo}���[�)S�HQQ�����ظ�=��q�����_i�s�|[��ͺJ�� �	F�1a�1c�Xx�XXɬ�l�S�Z=RQ��Sh�Y0i޼y2~�x�q�+�a,�z�@���@�!MK"��ŋ+���l(�����ٸCq��r��u>�A�H�,[���g�V/-.˗/���?''����͑��?_222$;{��5//W.����-�YY�V�H��u��6��q���0�4wh^�ȟ�|S,� 2k�]��!�h��Ha�X���%S
��92a���˼	ݒ�5$�+�����d��.�Ȯ#AY��-��)]})�ɲ2ڮ��!�m19X�i���ʧ���PC�m�P�e)%ʥ�ڥ�:Kꆲ�3 �guȎC��8r��䳋:ek�rNN�jж�������dDe�y�,�
D�d��9]��4G;V�� �O���7��w�ebn�O��AQ6��Wf��-�y�_(=��_5�i^��7���� �n��͚�I<7�-��5/	) ��7*������D�o0�T��֮���2�5uƴ^@�^������ֵ���j���?bm�,�IMkz�����ֲ�����BY��,�+�g�2AE�����o "5:n��As�m�%J�2��О.i^���K�!�5wiި�� d��r�[���G����$��:�|i�[�Uy^.ӦM��h����`��;Xnb��=���w���#2{�,9�:���z����c2w�\�l�1���*55��6�8ioo���F����ri--&����V˴^CC��1�YiM�Dӆ���Z9k@�2SJj2$�KU�QC�4Յ�E�ޑ#�U�d��)S���E����$Bt�$�W�ieD��r�.S��7��G#c��[��1�d����	F8�yn,�f�k���>��!uuu���ۍu#
��"E�¦(M�켌z�nkkS�5����ߔ�d�e�_6���@�2�eMM���!�������̥������˨G�C�����{ƟX]ce�G?<#��GOOOr<tW���ѣ&j}��-�&� #�7J�%�5Y����VF�CHk֬�ɓ'KGG����UV�Ze� Q ```@e|�TWW�$���.��@HXO^x�!�	�J�-2�����I�&Y�|�)}�0.ϔ1(�� ���\������A" ���!��7s����&�qS�  �{�����ߖ�+W�a\<�����e�]fk���\7j~D����I�OwK`�"��k�O	̍*!> �۹s�Mj0,�Hʜ
��ar��Ƃ $�c2��ȑ#f��t��2�ji�����Y�����7�'��(q�5sչ���ː��/c�y��qP���q*��Oo��:���3S1�ܦM�nEEE���jY�b����R�|�4�^s��F��!P�W�u:���L��
۷o��3eήd8��x�y��7�>�#C5P�@��:~�������p�|�W�Y+�Xc ,F���Ha�!��ӧ�5��HΘ,��Ҏ�"J }:^�X{z��6����+=�u�$ѥ����1ي �'��I��ի�c�b��Ա�y��Ek�_�D����3f���
���?6?�#e�	��C�i�o���}��GM����ʰ>J���/���۸��;�AE�����7��"9����p�O�[�t�\��+�y�����wݩH��}�{�$�.bq ���A~�ؘ������Ųt�4y�߶�u�_&ͪI�n���޸B^���5C}����?m��CG��l_������4�c�{���d���!�Z>K��@��v����Ȗm�r�Wj��2sz��9Y���۴ϕ�g����������{[+����Lfj�Jԉ���?6j$�%�s�=&b ����M,̜9S~������G��&s��G�'D��wݭm��&�QJ�ʯ�_v��u"5�Tt��%tx�������,�}�.,6N����Xd��=*��&���ϕ���R~4OV_|��4E��[6WJFd��OwTT���k��õJ�铤���RV���Jsg@�\8K�VFd����{��4��sR��}Α���[���5Wɡ}��}KYe��_����,+�!b�u��OJ�=v�%��ۏ�裏Ј�;�cJ�ӟ��a��_V�8 /���YF���Ɔz�U t�	n�K�n8�O�K��3S��ʄ��f���~e����}�����O��.��⠽�û����uލ�=���$��=	`"*r�z �y!=H�"��$�cP�"=���Fl��,Dy"���S�����-]�0�"LsLe�Ͽ�zx���G���:a���z	�7|\��immI*g�h�o��v.&�/��GB� �caڟ��C�yb{����3k�-��w�}��)���@�m�f��e �o|�V��q@O���$bS�'��S�k<��To�����C��M
�瞓/}�Kf����@☄^�nD�y���Q=��w1�aEbQ�j3��wl#���N3Y�.���@F����{fـ0��[o���r�k&e�@��{v�R|4)6|�,��yHߵh6��ON���|��&"`�c���φ����7�h����ȸ�~�/��3�! ��'HÄf.�f>�"R"C�B�;v���b���$wn�'i��L楗^2�v�ڵ��� �I���!��#����Sp�#�����r��9�%��O�ؒb�b�*����`����ȑ�!㤫���l~2�""��  Y����(u@\򤓉6'�A_n��;iw*.9U�.�z�	�|�<O�x�(y�q�7ʖ-[N@��Z[Z�M4A���:��T),��|2�7����(0��f������;ԏQ��tu�����7������%Ͼ�S-���7s[�bE@ڎ��!I�S���snIe�p�W�g֍�{6\�8�H��b�' ������N	+'�`ee�Y6tx:�6�������֜�C�u�2$��Y2�S���x������Y1ɻl����͔%�L5����������N����l�}(���l�aY҇��F�wR2�S)1!懄>��C�h��;s$��ݻ��S�?l���g�Z�H}�|[,Y�Rٻ���d�6�ʴ�C*͎��<5i�U��7���y�ޛ�`�&�2��D���@�H��	�aU(n�!�0Q�D\��[��l����w�+W^y���]w�e�qx'��P�٦��xA����ʖw�J���7�"l�|���Y5�ӓ�R�ψʄA����C�y������1\<:W����b�t��[�\����l��C�J���|g<�C-�9�ǽ��+���j�!N"�sVu���Ǩ���=�|O(��UY{�W_s��^u�������;,+�Н��e�ª�ќ3g�\�z�4V&�Iy��/��֓Ň#���y����!��I������APD��r��>����5����o���f`�Hxd�.����c�=&�<�ƫ���@�QW�R�u�� ������G�(�w��Gy��-���o}��ҧ�xB���ԔdKK�E @<2��k�Qjk�l�K�_�{A��X�Es�X�����"X���J��,J�p�ъF�<��~��%A��g,���k��`g#��<g͞=���m.? Jc�@�G-	0ʭ���$�p�"s��0�_� ��hl��Y3gK_o��< ��כܣ�@��nQ�l�Al F���l�ٛ�Қ:�d�x��a�A 2�|
�1X�w$?$�:�ebD�;� -�d�B/�����
"*�S:q�m O�`�'f{�j�q� ����=��s<^��,++I�8�)/�/���V&��cǪl;��K/M�E����6�S4�I&7� /K��l��Om����b�X4 eN��7z�Յ��b��aB��d��1@8�t:��Aux��
s
	d���|�:7���e�$�D����d�V�ѣUI3��VW�Z蜄N*Tj�8X����d��ܴ^������7����[o��a^�r�/_&6�ju�;������3�N�p�U��&�5B0�SI0`�.N|˙� �}�T��$�J����+s&���N�?��(2�Y��e�I"�W���_�w� ۷o�쉾���O����ig�%N��|��f�r���O`7�A[8F֬�cGsR%��C�$c8��C��������Ɔ���$���Mo��"���p���ş��v�|�o8�	����roy�Ώ�U�O�+�/��[p��c�:���t�=�q�ֹ ۴i֗�+_c�u��t=�&��0)��t/��(��S?]����yx���.� r��jY�l������-e�?���vp|���R�|�9���9���w���,��}���[! ?�;�ԁ\)�� yg�|�s��=���w�A�4�L֭��&WVv�8��1*�6�i�k�~J{�{gg�^�[�y��4I���7������:��ks��3��;��9pg�q�<:aTd+¹�x��K��͛7'�x4ł�,���<��}�D��L�l��T��$'�f�d�o�vB9�[�Α���H�����2�x�)�;���'p�w(���c�9�Q"��J=t�h�*F�4�/�d(���r8��d`s?��1 � y��ǒTw�Й&��c�G���N�>������ma���+�P��$Qq�vJ(yp1,
InR;�����c�vGd�Xsd�i�h82h�E� <�n�р=j
`38,Ɯ�����?�`�<|�� ')';C.��Hj��)ڧ�bF���F���a��uE�}���i���T퉠�E2<����pVcS�mK,�ܕ�P����'�|2����;aSz�D�I�&���9Ë&!68���IZ�z�W���k�R���&;'�޸�''�ᦨǲ\�x�NH�|ox�c~ZнW�7my�@��k֬U6�ׅ֞�)�/�~?�����s7�f�IvAzkk�9��p�4_=�u�]$-]�ޛN�ׇa��u1w�+e��.p�CF���ew36j;6H�_����P^8��s(�M*"�L������{v�A�+ s�z���D
[r�v4	J\�r��;�q,Z�0����+7�؉�R�� W8��)�Bq��8��<��.�8^x�tɈ7'KV�?_j�e4����z�'��)w��_������?��IC�"��X'NYpD�#6n��qԁ�	@�N9���Q���S��h#	MS�(5N%uu�I�F?9���5�u�p�D�� ��!� )~P���x�D��� [�.�-o�,8/6
��@wR�?��S�?�)ɞᐃ�w
;��q��h����'���������@� ��������㔢�%��+/�T� 0,�����\;�0<���{2��c1�`��	XZ���hYă��ڜ�FY�>V�,o���'M�'l�~���7���w�5'	������<��AO�cN��ku��w�<qB}��7��htPuG����U)zlR�q�=56wʿ?�S.��̓j9!��9έ�(�a^�Dc Ġ���)���n4J=pF�k�)���ݵk�\q�F�t�����5�\m�.Qx[�l=#�)�Pf͞m~D{{�����x��\���QnzY�1�LN��\�i�X[z��!���ALn�;���� ��p
F'5c ����j�(����Kd����M"䡇2d`��s��eQǘ$�w��i�=��W��&�1
��%8 44DT�u��2��	@���l�u��C�w��a1��@41�v9q��n�l$���W���XuHը8b��2�@�'�Һu��.;rq�%r��!���{F���2}/:g��ٽK�[�%��(CL�TU�*��Y�������"��&I{��ɣ�Wn�Z�C�xh�nG����{�X[��X����ok�-�h_]�6��i1����O�S����p�5:{��g��?��-�@)sWJ:��/���"�1���{���;� i��-v�=��E�{����?�)�o��¡?�@�D��?����K�ͪ�I�wt���XnW1�.1��a�bU1�_��I����nR�q�!fӦM����&ĭXڀ��F�|o��G�\�`!�`�V+{�|b'T�9D��ܹ˨������O�: ]$����Q��7s�-��C� <��g����X��Sb�.��q���+A7����o$�d��#1���o��V�����0�pi�3�''���	����GW	�p�ȯ�s<�& jZ�����͕g�:��񹤧�F�?%B��v,@�'�}h(�Is_�|D�}���ZX��@"J�;(??��=�#����T�`�|��7n�h��������0�&��S�T�2���|��=	 �D�'��]P�AL�Y�s`<8D�!�p�� �."}BC�����{��6��k���g��!?�я��1 ��<|���;����H8�{��N��wؠ ����C�	���loo_�T��t�b@�7ސ@x�!��U�M�v�r PW�(����%�䉿| �a�46u��ͫ�6|"3�Ȣ�)��3[e��n�:<$�^�(��fI��,������_]-7�ܜ-�-xz�����-�o�{���������3�d��VG�to����er��.�Y�Չ�hė���n��6�Ǯ|�~��X�'�0�GM�{':�`g�> �/��5�T����-�
k$ l���u���޶mۓN�By��]��;�j��˃m��m��?����v�0a����N�R���Aff�|�����I�1�m����6$/m|��|����[�hlD�}`����+)���7�R��ȯެ\�f�������]}I1�KB-���C�9�湚�Y�pe��w���I� �.��rS��^{�Ev����N��'f�肛� Āg�t�����17n�`�n��H�\gN��R�!�T�}��_���&ikm��7�r��|RbD�q7�Ζ- CgaX@$lJ���{���믿a��H�K,S7|85ÁA��f ��LD�2��/7
�W�O2q}�w�S��$���<ŷ��~I�fͅ#a.  ��t��������"���I���Y ���=�nx�׌��N �{LZ���C���m|%"8>4(�� �4��-��Q��}��Z��BԀgNUr��q;:��q%��z@
Ҁ�p�K��bg{��PX/D����`�:͉mO�7�e��!�X���apFA<���i�����|�t�Ꙥ�$��&
�6l�`�P���2Bh��X< g�hD%��m0�$��@,�F�S��v?��~B�2 J=?�ȸ����pm���[%�M�Dz&�OK�i�)�!�Q� M��� 0�{Vv�����^�ó�se�v�.#3؛��갽DA4=���������fZ��tE���s����mjb$Q���`���)ត_���Civ�`p��ʘ�#,ħ���Iܔ�b�'M�K;��_����7]���\�!-�
M�ć�-ґ�"P*E��@r�R͗i~-T�u�	!�˦Ș��-c2��`}��� ���.��L+��]j*��R?d���E�T$�`N�1߄�y:����w��<3/N��V������A9gZ�mJ�±�"��i]Rѐ)�pf���Z<�[��f�$E�}K�xj���4D����H�J��dQ��>)��+%U�F ��̊�ɬ��R�e
e9�2�`@ʪ3�:��e�ȸ�9P�mđ@�?h��|#�z���B�@�����%�e��2�d�G�C��=h�
�b���w�xW�e�ǝ-��3h���dN4��Bz�^c����ײ�.��� ^`�O�뗺6��z�(`R��}u��?��`Pv�N���}q�?)�_��)���nv4��U�%����hB��/�ٸ%��\f,.�$^���o������˅�g5�)�� ��H�{;��[%�#���+�C|Hٴ1���Xd��c�x_m �"i�Z�d��Tei��F+�q$7�>-k��my|bQz���ݨ���|s���Ղ�z��/��ޮd�|���̞�;]�\�(+0�tuv$O��QVh�X�x��_�h�-��.I����Ҏ�F����2�^��ʽ�3[�;��Nb�* ʫ[���%���9�DZ�Ȩ��D>�?��M3����/g����PrX;��B^��4r�= KBibY��~V�&|���o"��!\�s�X,�CY�.�@�a�����n�����8��Q�E�B&��_%�9���O-R�a����e ��y��2��_q�Oq� d@����������    IEND�B`�PK   �eX� ��! �3 /   images/adef7304-bf01-4449-bba8-564470ca0600.pngd{eP\A��������݃���u��%�BBܝ �%�Kp�`����߭�����vg��������5�1���@ ����.��!��B�	���TwC/(���.��^�%�����7[o?O����������������	2��� ���a�A1��T=o!�Ŗٖ���A���GT噧cԅr�k��,����vH58Q�ͤq�������Å3x�HI^c�P�~Q{��gxei{�v�Jv�"�����pI��í�m��͔	��8�g� ��v)�Ep+uc�aʪ�b	D���� O��8x��A������#�֟���OQ<#�����F�[�<Q�kU_,j	����},��php��E�l�z���:^)�����z�o�FR"��:���y���B�	��.���'�җ9����l�휗9d	>��z�w�/s��#�Ү?��@��C�]��s9�����D�z>�RF!�Xj��h�G��rѩg[xq�h��2�i�����$id&�`EQ��R,楚�Pĩ�W^ }��ƽ܅c��??���`.q���d���/*�
�9S���L�(���{���8��j��ѹ���b��Mҥ�����U��#I���ջlA���G�,��ϐH)l��̑�������Ļ����Ĳ!��jV�H��`bG�ϻ�2.q�",̮����H���r��1#��OVp5�-A�[��%��q���H��]���<9�6��&EB�(R���n"0��_�մ�9Z	b�@���&�ghk����������.n��x�}Z�V����!���UT8���<<
]�`����s�ǔ���{��x:_�7�K�!���B��Q:9ځ�)��+Gг����蒖t��d�E+�^4j-���?�|b઺=hzQ�w��)!�nա�9��
�-�W�_kVg��Qe��7et�R����edע�g���T��{T�q�O/dՐ>�o����5c�,�����}xW�$x�)o��_���ƈ�8�2�z�#��7~hP��4�h��}�/���'z������و��ޟ^r���}pCY�E��~� �p�J���Q��[�y�f��� q�+FO)#�$���9)�Y�����������o�*�*�����]�{�3���Ji�<�e�y:ɣ{��U4�bf��߮	͛ͮ��e�i�<�#����~g��Ro(�8�EA�{�`��A�������ټ6JńY�-+��+��ȤX��o֚˙���6�J��}�	�`B>B:�_uI*	�����VB_@�q��������r�����l�����7�t�<�D�ë�uD�Hw��jjǢCS����t�H[`}KL�O�38����݇���R@AzE�h�"��n�T��Iy�.���.���^y
?ܲ��f�;�i�3SU�N�Ä��	��{J��� �z�@�������[s}{]�,�i+E`ЙV�:�y����ïH��wy{)N�o;���^<l�~Ic�
�������w�Z=%�^�X	�ů���NWD
�j�d<�N-ۮl�
{E��������|����=���?}�"�$� ��#���(�vG"����
��P��?D�zr ��j���`�����l��0e�z}�~X��q��S�i�Qʸ���A��a%�;>�l�5EG`���ul$��̍#�EOC5�G�>}�Br�0��8�"=L�o�]x'�^���wxz��~�S���.��NA�d���Z�p�~4��Y-Ƕ��=�L��q�̸WO�s�*{���Qf�)%��H�¤��:���� �K25��eË�%y��@q���	K�"�ŗ�c�/���4���oxY�[�	ت���"}?>�eF2��(*8�@&	|���%/��b��$�m�
@V"�83�`Q�������c��D��Fx^,g�WeN�R^M6Ŷl �j&O�DE�^���� ʍ�G����s��Ʋq��r��xVa�*x=�^�pEt}��҂���k�$/�� �K+��v?I��$iߞU�M���2�;�;q�1��b$��a�,��[څ�f[c�Q��Ř�(�c�����ڲw!&/c�3�������Tm�㉗����nW��7����-��r瓚'!�`B���
���>Pb�a!�������M���p���u/pz��Ӵ�s�'L&2�&�R�MY?� ���B�֞>/̂+�]�����`�R<va�LZȟi�*i=���)z����ē1|Y�D�"�QA =�3�`�2�b-�����r�/Y-	G��tk+h����^&Z�b3�I��/�M�@}uf/�ሺ��:�b�Y��x����ǳ��զۭ�^`��<II�L<�ۖ@��z>wD�:I$1((��{������}7�.6鯿��XdYX��J�;���h����0�1LO�78
�����������5u	T-���?�œ���Z����Ya:r%��<��W�S���i��e�0�s9�hi��I�)���OU��t�u���6x���zA���}��l����d	�1��ˀ��7��^����S?�ʺk��O�bG�����3{����⬰�pQ��Z��'�7�s����J���=������m����$�Nrca��Bn����٦4�cЅ�(�nTTACz�� bg�ϠU)�n�2�g�kƹ$��_�ߠM͞��T�u��R}>!�s�U:��9�����y�QQtLEc�wT+,����W��s�7��4v%:#JmiD�ٕr�2��S˲$�U���E����5�C�e+2���B�&��P�?8q�ʘk�`�0m&9����9Ë�Zﬀe'P{Џ>�N~y�aܑ�,���h�>��cY��E-�D�x�'�Нv�O	�T�u-Q ��$�(Q�4-ZI��ړKI�J�ײ��Jr���.j�Z�L�#~%�J�s��&fEyq��yjB��?rO}�i2��������Fz��_o��(ŠId2;�P����q��@�Z2&�ؓj�F�^	s-��u���^ �xG.?��d�5���W��+�|��-�^�%{92'��z���K]V��O{ou1�N� *�,
�0~Ca�(%�?��-fx��*�b�= ��i�<M��Kc�z�J��b�'���Mw�d�3�*@�&G�_��*jW\�:�W�z�"��hF&�--�^�6:p�S������ͫ�N։��KL����L���e�R���2�� �GǸKǵ�^�^ u�H���EJ�#�����V*�	�g�m�����9���"\-���%��d�/���#�F#ˋ[6����t秫�wf�ӮTF�ߟ���+�G����H�`�mW�9�X+:�K�25풮���_���8�a�
&�G0�Ac��.hP5�_X�Y���b��]��0�޳	�K�#a�54K'�
 ǂj-F�}�z�
�totIo�/y����b��5��!�h��T��D�������N�݌�r����ԛYOʸRnIJ�ym�-���g�:�n�I��.WU6E���;m������6����T=Wb1igG�ԍ�~�h�8���}�����D+	�#���Z3	�w͒��U�^Hc ?�jn��p ��|#������% d7$�Ю*ǝ��4\)V?TP��PbW�mN<���'ؑH�ZbջH��,�i�����!�����]���� �c�3*��Z���tG���pؐ33dS��Tу���1��s~�>fd���+�	����_�ӓc��?�.���b��УA��;+�����I���J<��am'La�l��������;���dͶ�!u���
x�]��=sSq�UVi�Qb_�M3��Fv��t�6�J�Fv-���fki�B�('�Y�FJà��s�kiW���P[�p?4		�Y9��.������֙x>>V1�0`���TNLSd��y�0����!��#�v0��E��%<TK��,C��z$�6�}�����V��A
W���y��P���������W�G�2'r������Я!�Xǎb���o�Wﻈ��1FZWi�\�Q��_Κ��JFQ�{�׻�:Q�܋�>�?ny�"*�U��#��?��r�FJ7Q�D6z��5���()��E*��708�J�}?	�`:�O�4�4}��1�� �F����]�@�Lͣ�L��ۊh�����|��F�4��ݥ�����O-����-��誰��!��vOr;͇���1�0�o� -:�l��\d!���+'֗O)���wͰ$�L�S��Z�,��/`���@��{�@@bA���9]��q� ����Bˁ�7UeݭQ�YG���s��=�J������GN�w.�E%/���v��/����hʡ[�"Ek՞����Nt�`�
D�������H!�GO����S�	;�UP��t8b� cL�A�=MG���' ��T��-KH��KG���:)e3Y����������Xw��mĆ�����x~�����<���l����M�}��\�`�i+��M�gzu�]�ՀA<��Ԣ���O��4L��⏢����cɋ��7�$_%���W�
��n~Jh�/:H����|�')7?���'@�|JR侄)L;����R隭�����0�/��n���W�E�ܢ��&�E���{�Oo��|d��MM��'����\���c�H�#�c���?<�2�Ua(���}^��"����>֫�����U�k�nK��l&�K�ۏ�F�2�fc��$Ǿi@}�c܇��.��)��I᥃��И�a�s�-������ƿ0���9��ó��_7e �rſ���!����U� Ds0E��X)e��i���-�8�b��O�؅~�1"Be%ݼlD�\^��|�4��E#���є��uV��"f�_da>���3�!�8������|D��_;l�"Ҟ|�>{z��m����I���i#�(Mx=�5��рA�Dq��?����7�y~.��C�����!�j�q=]O~��^�}��-�L��eaI ��.����{��sH}aB~"�r(t��=fW��u}�z�{f����t�΀F��r�ZHWtB>s�i��#�b~�L,z3ܶ�|31Y'�x�k�:m͕Niɩ��)�f������O�3��o���I�"T[�J$���~U�oh�B\�Vx���X�����LK�����T���'���V�o]���܂�ECM0-zS�d��EM��c��â��n�U�A���]�J�w�sg�C�}��P$l��:�n������U^Z��P���&���o�-��w�6���W�Y�Z����|�jU<W�|r��:,�B8!vcբ�v�#�		�d�a���)pۢ��񟔡�_1B�&~���e�shF��.�®+��!|B�y������R����/4�L~Ws�fЅY=��3x�/��t������߇@_��kv���{�����@X�˟|���H��1����
w��#��ݼ1f���Đ�dv|i��47%x�������A���a�=�K�E��\���Y�?�m»��A��ju��Y�eD�vE�~���&�1�ްXڏ{�s�tD�y�ῗu�mK-z��廪��ɛ���L���2�fd���Zb=3^J�!����Lzc����#���	C@�B:��η�Z#q6�T\Z����M�f�Z��υ��nd#YX�$�󀾣��V1Moa�<PB.o��^����%T^�ڣ�JVSmC��P4�*��󒿌�^9A��Jbw^�6�滚����]��M������4��A��S�y�)��.�����j�+֌�2M��*L���X��_K�|&;�^V<��,�~cͻ^�}�߇����53��P�ճ�Ɩ�E;�8����Sr�KJX�\����.-g����i�4��Tp�"��@�M��)K��mR��(���I�>��]ރ7��?z�>8T��a�N}~���HU�Jh�WX�a��LV�C�-Q+&w���x\����[��b���=|nu[IFӒ�����g�q|/�n��G�^�	X<|�b��o�w��n�'��8llC�h�����I�� #�Q���`�����Ev�y�̫�=��v~uRBu�-\z�$�zf'!�ی�KP?rZ�J�앯�w���k����yH��'��K��Eќ�G�H����@'��#&�����'�R�.��Lb��(1���)79�aq�!d���`!�m��<��S�ו5�dO-�E��\��P��4:��O~e��^�͏�Z����x�pW�]��p���B	������-�%V�*�z���w�����iiy��{�Q�'�c'*���W`2F~�w�]s��`��? ��8��+���#����~GԷ�L����fm�ݝ�e���C�[��4�_�����0/�Fxu�<j�������Tw�Rf^��i`4f$ ʎ)��px�CNW�)�'����"6� Y�� �P~�,�,����Ik|���I�0]�5 ��҈��t�d�d��m���<�q���C9�k&���;v��K
�Di��	o��Ĕ�;"t�̥��߆��`D6�GB�R��g#?���0-���%M���c����8N�+I���FH�8��M���QGr��1�9���M&4�|��<1\Ƴ��S?};�(T�QRմ��������Kj�<UT��w.9��Ƃ��W]|s���մ�`�ѣ�ܨ��IB�}o9��}+wa ���)A&e"��S�f]^}ɸ�'�i����kw��4��Sek�L\�_1W6t�Bo��_E�X���~'����=���>d��$�C����т��uj?�KOԬw��Q=�I�H�)����4��k�Snc?����0W:)D�Us����.���T���L�Ј��א_�`�x�9U��*��?ކ�n'xe.�H��IbG�bV�Y��bw%2�`ǝ1�F�ڷ�����QKV�
{xd���ț���Z�<���\5�����oY�\RWry���J�UT �5���X�EE�	�ӫ ��C��d�� v�?�k�%T�bu�����ܪ�� ��*E�4��ߑ�]�dIPۥ_N��X�񸓼�n8��6��7�K�j[�G�B�]T�W��N:�}�[�*�1�;����Y3�;��.�Ru뀟�"��~-3:�ug<��g�L�#�I������r�C��"�<�z'��뙼�ET�(g�hP;\�8�q�͵��9 �%!�Y�O�����W�I�0+�"C�v���]�K[KLܽY�h	ie� ejf�He��������[�C��]E�� �99�>#ۍ\���tq��fW�#�������p;�[?蟓XmA;F����awjM��w�A���+t��!���Y���nץnt�!�1�b7U��c��.��<պy6�)��3�giQ
���T���+��k���J�v� ��[���Iǌ���!�N{���zQV��%L��^������@�t����|1��� ~a�}u�)��1nt=��2�#��N���6�9������Q�IDK��\��������Pǭt�η��}��v$�_�[^v�bFKk�Ƹ($���ͧ��e�'�6�x_��9�F�ږ���,/IBI;�lQB�N>@�U�ȟn�i	il�mOL���#u.��[�^����:��$!���^�q�䭭Er@U�P�+fʡ�/��Ao5Y���	2�����p�Y8
c�#ؼ}�h֙�bH&�p��ޢ-���O-Ufs�G���-{�8�M���c}"T�d���} 6V���M��u��H���Y�=13~�����*�Qyu�v.���Կˋ���T����D�����C�ώ��ꂴR���>���c��]7/�e��9��L�g�
Z��1�h$�q���V}1�60f���I�ۃ�=37}����E�vtT�W��Lj[�HY6��f�cG��f��=x$H�La��ub����.���y�FLR�|�N-=��v��_T~?q'��9GnJT�޲}��D$��m�rb������v3149�(w��ܩiyV������Y��P���)��RĮ��*V��[��_7i���8E揷�ڦ��$���(�@{l�"Z�]�#_'9�lO�o�cж�T������gs�)�LH<ұ�����g�����"X�,��Z���E������|��ղK��0�}	�17^�z���mVq�!��?]��W��2�rhT��Ր#�`W6��TX�Ҧ��mZ��ƅ���cn��Վ�<��O���r�|-��,[�,
6Hˠ
�#�|HN�w��W����(>�-H��{��c�%L~(�+��J+��r��96+(�	���hל6ͪp�H�{��{�8��E��B\_(����t�*{n�6�ݫ���
91˵7�Z���E�6����ܦ�?g��՞��j���PY]�~��_@��囬���̒�<M�{D5��{����J���[� �!��7��񛔏�c�ba��}N�)�����j�G鶬�1S�٬L�a�%Ҙ�Ť����\)@����4��������lV؍��m� �E�"9/�K��b�eC��K�qw�t��}$�W����g��{�����;����x_��'kf}�u��e����1�U�篆�k�7�|<�+j</�I)����P>d\�����	����ڧ4Eq�xvW���l�t(�z�:�H��=j����Nf̉��F�F��͇��o�!C��q�" �'�����4�5�[S����w+)�=o�ܔZ;
�9�Y�Q���G3����W��a�PV�	�@%�z- ����&¾�gb���*g�i�'���$#�i����_�J�|�u�;��r;�T��G�q�u!p[���v0���ܴo�%5�8P�L! f�k��z)|���o4c��c?YP
^����M�EHg7�o�07y_���2Ƕ��Lj�w�S��m�0�_�Xk��DǴ+��v�
���m�KO�<S����U�_�o�3i�FP2eO"\絴Ay���0���4�86y��QW3	���J�s�zY�����8*TX�������0=MG����(��(#R�q����a,���(��۞�}�0��6�wC�ߖ��0�F[���(��ٹ����b�'���j�[�y��k>���Q5��mqVE)��:!sC�[�3ʸ�_�4u��K������(�C���`j�V�
�����J�4�������<~�O뾋�cl�v�Xt�N���~Rn?���`�
�RjHV%Mu�+"�2�����d�K�r�eF�)A����nL�5d6��q���m��ʿ`:����N�g@Q�nqF��J��}2,�-p���F�.�t����^�@B�����A3(�������j�6���@��v��#�Ƚ1�T��P�J�q�a�	Rh@�k!��mNR��*�V���Ns#�;5T�K��Fd����b`>]٨(��5��T�*����;���Դ��.�V������:����#����vO�1C�M͗���1�%R_�O"q��;(G�J�5���c�y�1
"�ԑ�K3���]"�F��1��gM�f����E����[^[������xݾ�z]4�n��������enNB�>'!���KԢ3��n�5v��#~�L��aJ��������R���5�[�^��Ư#yJ%փ��[���=[9
��;�i&���赏(��>p��,�]vV(����DV�kC_w]&�!��.p�8��8`��-Q��vũA<⢨Ǻ����o�m����=�?�~f��2o�+Ĳ5�ب>��`*K��~��X���m;�ʷ��n��Ն�6w̩���a���&e(�~��s���KWf��0��ϧ�RK&�2�i!�zڊ�ay�H���\�R5k�Tc���Ц^	",�,�h<�0�7�����}�~/���Z��H&)��5�IY�
��� �hDY�F�E� ��;�m��`1��⌳%�i���o4}x~�Ti�2.�)D/�]�U"��(8 -�}�\5v���i������:�80�,Z����	�+oXJ�Rs'$�;$?BE�i��y\�ZL���ۿ�������sn%9>�^����p���kt�����M��'�₳���T:�~R�Jz`'$ŏ/����S�	�9���=�{*a��+Sd2���S�Bbmc�q�	�/���*����k�x5��%_V�>Ӱ/-�n��#�ɠ�R�W�6�����23�9�l���N�e}x���E�˱\�,��K]����YG!Ʀ��آ
S�xu�H�-Ȫ*�!7�L�����^��
��xS���PEl�Di�
�L$v�N@���592���$%EKEIדi nxC�pϯG�~U0�)�"�me뫪���T�2=F^|������Pl�������)$�^�!68XL���!]���N}\�j����"���0qb��T��K";�?�����E��Q�l��DĲ'�pމ���v�*zH�n�R8k���n.e����%3O�(��]�K$�8���`���@��X�嘯���=v(�44��3�<�q6��?���]�:�M�����#�(�_q��0"�p\����+Q׷h)�"�
Jf�Dr�B���J�Q����x]2U�zUO5��s�
���v�̣6��m��5%>�BA�m�ه0�*�pe��e4-Ҥ���RW�U?�DN�F*:U$󎜠��(�?aj/rG��dۊ���)�Ψ,w'D��;��Kga�i_/K'Vx�A̪R�����9��J8���Cj�]�^����|q|�����N��5�}�&@/�M�"M�>Y���]�Z�
�V�ZU�A��u䔖w$�$sS虳'�/C@�s-�ȣ0p�Ԋ�H�6�q��ǩI 6���QW���"�	r;�}�9�ϰ����(V[�YG�RZ�K|���%~?Ib����@�*M���㊭�3�iz�]"��:V�q\J�����al�t:|>�8��V��A�u��<�$�q����@ۺ�
��9����ީڈ֐��OQ�~&����?!Kۛ�0zg�)�n����`�Oa��
��n�O��}��B�?6c��G�8���1�}@������!�9E�e����|�4
$ݲY��j�D��I��@��K:ڱ��0�5?F�}|�����#�k�a �p��x�;d�z�<Qf�O;J�| Qj�
n�=�kOj��.���[8Yr���(��3��&L��Я�_�_t���T��L>�rR��'���ӫ�몢�4`>Ja/�GuI�A����B�S��!
��!2wK��%�,!q�ag�)e.������׆@�}չ�T�nY�a����7��oUVGl�ӱr>^�T:���O��8=/� �78�{׏P���:�^i�K��u�`޼�*[�*�����t6x��d��\�WQ��0��x4TB�C�P��[*�Ph0�_���o�g�@4NE��*�:!��6�=pVLp;�����i#9�!RB���!�a�lx�g��Hf���J¹�8����L�e�ƨ���i�D�$��gQ��r� b/\�8b�-��)�.�!Yޑb�~�Do����3��?�Qhّ� �' �a�t$l-���-��HB�R��T��*'�p,�^�]��Θt:��-B�rroMd���s�rãx'�~F���`�S�"��͠���)#L�?%�!��E�E��Y@�)�<��m�-:���>E�z���̩�N#���A�ސ\X�-�KBTga#$���V�����f3���Sd64}�v�k
�29�QSҢi��e�:z��B惛���ՔOi��

Csl��9XI\-��̧N���e��1�-�oZ����A�Td���7�+��0zYn�/c���&�48g%M�X����jԄ���=ƱR��d���ypS��zHd���+r��Ƒ�̏��|fƍ}�du�~}c���&q�sZO���G���7
���S#t'�:�ہ<ǡ���-�f����8�!�	x�\H�<��0U$Y[���8�k&��z����գnY��R��n�f�Kjv��wh����b���֏����(��/0[PB�)���%>��i|j��BJ�k�sM͹���v����Nj�s�/��68�b��*ѱ�!L���Bt�}iZ��n���J�W����v�|��㏁���K�"E�M�LT�5**��������]����;<yVC�!�����7�;�@&'�v��s �U�7���9�EI'Vj
+!HUYZ_�$���/��:��`���[�~�MU��U��K���f�e��vO�!S��/�N��6܋s2���X�z�:���͚��3e�':�2)��My�y�<31�� x�N��g>�5�5�v&��_c���0n����4���4?i��L�L@��\���	`O+̙��H����B� !��m2ݱ߈Ǧx]��X�Ô��QA8Xd�d��g��w#���޾(Z�IP'��ܕ�Y��՞cv
�A�yq\���
� �wb��=�L�I��y� ֩��e�� ����
A�3r���"��S��j���
�����W�9%B���^Y�鵏�Sq�HHO�����Zx�Z��C��I���D �͈E_l�S=�=Sx�>cp��|�h�®�D[�=9!K8]Y�F�� I�-M����\u��8�h�wЯ��B�|���ɭ���D�ˉ@ 
�3f�����1(mO@�ĥ�����ئ��@q0����E`1���T���L��qK��`\��/}���^n�` ���i��8BO�9��Ht���m��%^�^ݍ���j,"�	�+�C1�� ��~4���J����D��Rrʋ�{XM8(�f��|W��X<�ߎ�N�J>��R^"d�rn�n��;3��(ʞ�Cy�K2�Z7�I ���#�c�L�g`��#�kݽ}�`o����#�G\)Ξ���"�������'� �j�G���S�_P�#����.q<Z���џ�Z���dȰ9�	��n.�k��w�%�sYn�~�-Xrs��j�M����e��A&�Q��1f�M?�=�J�� p)��9���IV(�b�J/?�mŮ�J�6�iҒY�g^��	�/:z�;{g�74���æ�q��ӼtY��4��hϭaI�1��řD;w����?��a,۷�V�,�ݞ:�;�q4�T/}�X���Q�+`?�QgdoJ ����_�Y��>/স�Ce��iդ�����0��n΍i���ز��m�*�UQ����q('[����|Ӄ�f��L>��]�J,��3I���S��fN4�Q�<M�A��[���V�����L^|��� M~-˩b�6�`�ɾk��R
9VE����a�9�,s:���H29ֶvP���0>���ۮ+�s���;�ͳ��]�Ԋx6�<_Ƥf�
���-��eu֊%������?�A\j۷_��K���D2��W��.�5a��%EII�]���	�u��l����xO�{�|�KM���ۤ��A�>V����h؄Գ��Q�r��uq���`�n����]�g���_G����������<5��ޑ3	�(��o��G���(�uS9� �����v���iY.f�C�Z��z��h�=��4�/!|$Y|�\1�l_�+!��I�lp���]j� U,���E<z��y�P���}c_��Xo��"��R��"Ķ~���,}�J�ː�k�nl��f	7����-E6mN)P������$ F�(L*v�T���w���0g�[/��U�E��h\�y؟R�Ս*w�T��������};+zF��<���JBMޛ|S;5���f򥟈CFnCH�)8؋	\��&X8k� Bk���l�ec5�{�r���{Qek�hf��-!҃t %1,9/�ڈ�{}�6T�!I���JxY�C�����>�����ֱ�sts�遌
�H�c�5���I6�c���G*t�lRՀ����q1�d��*�:���ⱈwG�2�ȯ��D&��Bs��Ӷ� @��E�����\�?�F��w���qNN�R��>��F5ل��<�|8�Ve�fHK�1�:Ǵ�X��"j��y�����B�k��&���_�(�xAE�,��NC�䞫02��|w3�;�Zg"�Ժ��kQ� 8���xA���J��=�O���Ob�zst�2���4<�ӧ�v�VH��3E듫¸���&����=���[S���f��an�-��We"|0�6S��'k��oJ!}E�I�$3w/�Ŵ���t�a�;U�?��Y/c"���4�N��op[��~^�s[�����n�8D�)�mNߍ)�9:X��Y�Q0kC9[MT��f�*���;�joUTQ����W�X���8p��'0�$˫%�d	R_��<��6��c��\)�l�I3gn�(tf��!
��j�jI��(�~��4���]����S�)�"WZak�a�|�����Uv���'������c�(�CKNP�/�[�;��ə�5�@i�Y��'�F�{]�7Y���l��������\I����!�N�L(��̥l!ϫZ�W���;�@K#L����7]k\�2Q��$�y��sZ �ȅ��Ϲೃ�Kk������ҊSk���c*qa�U�j9n��ϖ��=P�u��b~5�[�@+X��|�|ۡm� qx�r�e;�<��������o	�+�:1Ӽ�ӝ��MS`]ڹ|�u��FB��+��)���7�C)�����q�K͵17?��X�I����[����䭣���]L��k+��M�'Hf��"���Yq���Y��/�6q.�����E�*;K�LJ���߸�x�o��u[8���<X�*{��H��J�.����=wq�7Ҫm���h�Q�(`���k�@n��i{5�n\����[�Kfa7lg� �MVU�L�ʺP#ޫ~xz����e:�����)��w�f�Xd�{�֍C�߆6��i9�-I�te�fl��� ���0��G1����A�L��H~�0�V7��޽a��G�s�Z?��Js�	�i:0�&\�{�~s�i���d'���ī�m���?�2�8���K����O,B����q�)K�|�Dv����Vsd�w�"���]�u�26u$iO�,�y*p����n�݈�b/���p�ݛ��µҎ5�Q�d��V4��D���b;�9�E��痤נM|]9@:V�E>��S,>�x�	��&]���C��8�dǑ���|P��`+?@�1��S�Ԑ���`۳�6��/�����wQ�5B�p�-T�q�;â��d����yս؂Ui$�)V(1A}4=����.�,{���t�ƭ����%�Н��g	~�L��	��+�^�9�ןo.p1��@C�*�b$��ς��B;�ՙt��7�G�G�ϭb���/����3����z���@�&��\���"��"/`*Q��Dy�]�艐�·�M-u.c1���ԁY���v��P��0��	�ID�j��SD���	��zy����
JY�!�v�#$��֝;�5�Gb�~V�{�����,�{w�s�].��>M}�e|]I�h�\���i��9{ ����-���!S�g����'}Er@�^��*6௯)� �vO�/��S��S����d,s�bt �&yc�hH&$�h�,��t�=���R�y{���f%�m�fh����=k�z�wH�W�F�@�w�,����/J]0�۩��GP���*,R�Ϗ�G��I�����9�`,��Ѓ��E��Ϥĳy�gn�؏���+³{��T��޹#b?�� K1Ж��.!����|7Ϙ598�[r9�yU�꺁�џ�54�L���݇u�I۱�<	n�6DR$5X=.�>��� �4�Au��懎|��V�+.�s��6t�D��,�p�@��C2�bj�C@��(����`����y Y1���eim_g&&0��w*V鞐�?���_Y��QsZ6��|�T��u��_3�_�K]x�G$�g6�8g��몎ݯ�#�J|�.̯�Ԕ�&������X��cn�'[�G��J�N���J[6���_�$Lo�>1�J�;���[�/�$��ZL5��
�O�,��RP�+�s��y���y���9z�lVr�G)O�T;�B��%BOM"O�n���N6V㈮��d��&�k[b`d�����ǳ�v��B��Y[��5՟Ȑ�ˉR�2�E��U}d��	�8@	i����2��B�N[I���=a���$���S���.�W_������b��jֈsb�]_]����f�s�Ur�dr=����³S�k`D�\~B���Y	����Hǜ	ъ���aL�s���#-褕�k��%H�Խ&%��I���#�K�
U;t��Ŝu��*5�<N��r+D$C=�������y���z?�#dP)Μq�K���J�8��n��ə�N�4�������5�5Ì䉏 8ž���n�o���ܕ�	6R���� ����~|	��C)š:~�����5��Uۭ&QqZ}���8#k�;0�H��������C*�ﲾ�CfQ�vkC����"�gY�����[�E���CI�� "  �4�"��"��(% !�]R���H�8�H=�5���;�}�s}����y��b��^�Y�z���g��'���0��f���:w�tg$�	fV��?8�q^p�/^�f�ym�!����/K�h����-�*���^]�l�q>�Rܲ�����a�I�¡|dKT����������)GQ�'Z�X�
�aY5��Y���QV(}˝�{�5)#�	���k����E������O΅ì,V��F���	[^<�[=͒a��ǜ�x}�O>��̞���}�y+���_i���� xI�8�Of^�=��R�#����ƛ��G�9dD�7`��z�4��8�3P�!�Nxވ��/R�>S����+$�� �.ġo?<�W%	ݘ؝�~|�q~*f������p�Ʊ�Js�M�s�4��W��\�+7B��xc��婙���3J1�����=ϩ<��͍��,�!
M)�'-���}���zu�9�?*�q�x_��D�.�R�A.-7�$��F�]�CU�� ��j�&B�C�ӓ@0J7P�=�+y�M�����I�گ��>5������sx���������;տ\-�"@�k]&�^���!W��Aa]��F*�]O��T�����:�����ٓ�����k��4�}�
�r�r�zT�G��/�d�����WO�i���~��|�<�v�l�?�-����w+�i�]�=^�Y�Ԕ؂`��_��_�<�<���Kq�����>�dm���h�C!�u��/6���gM�Y������`��������}�*G�.�|��~&��u?�MG�R�����J��#x�z��+kF���k(E��<o���_�:��x�智�e��ҋ�����������i�N��g��.�p4|����g�C8y��m��k\��oK���wAB�<�Ql���׻h�3
�����f�3I\�����DLǌc&���:�>7i����	�O>�i��9q�A��Z��m�j��ǴRѶ�$M�>��7�'\�V�4sW�-��!.Fx�.B3g/���~��d��[��!���9�cZE��:RC��8�o?~ӽ�����s��g8��C�[�2�4V'����u�i��.�\)��L7;±!3J�>�jU&��^��=$i��Lw5�_��;����qr��s#u��]�m���"��U����^�_�mb.P����������+Gh�;�%�L���Iy�^Ȉ�v�<�Bh����~����諴\�y���܇��a(*nrc"i+���2N����mځ�	��;���q��^�i5G	ߖ����i�A0����1�������;�>�^^<���G��x�
6kZn6����E�}^����H�P�>r�@f�
;D�gԕ�9�>�dL��#Q�xN���h���W�%e2[�'�>,�g,��
J;�ӘG��?}r�N��0�AR@�Pa"����)�)���/�*ve�P���2w]�>ؙ���]4�M�}y��?�e�W��{���$�9^�8+P58Ny�>��8�j�t������s��JR��I[�����E�w�^��DA�`�v��p��Nwb2��P�����?I��=�ťxwf�}����eTA^�T�7������q���33����x�Y2�� +��-V�aՇ$_p~*5�e���uw4p~~�_v� 3d��B�pPk�%�\��T�<����yL�0�J���]�L,��zDH�ʚN�`�'�G�Jc���IF��3���x2�+�l�`#�~P����U�E�'_OeT��O��A��ʬ@1����A~�'�I�f
!�n!Wt:w�c�|7��3�!�+
�z(sRH��sS�>~Od����x��d�����su����\�/��f,)�ψŉ�H�*��o�u2l����������Ē����u�x�9xe^_Z�W<#�S>�{�G�7`�_f3��ə1�+_��b�]�7������~��L����`�9��[x��Fő`���ٸ�I"W�p!�gx�Q��=�Bd�~�퍻����|�t�,��G��fV:+��*}�U�=?�!�<�	l՛����BaQ���H�Wrи�bd�<e��ٰ�>d�Pr�q���}JdΣ�w���D��C�q������z�~������.?�x�<U��[�W3|6W�RCX>+8�I�ֳ���b��Bw�^�$�Ѯ�t���7yQ����������*��1�5x72
����v��w��;SN3����}R�*]�Е�ӳ���+z2g����E������׫(�`�kg���+�"���0u��%ٺ�u[Qˡ��ʳ0*���j���_�A��'�|_�~�1x�Z����R���U��|`��>u�Z8J2�񙸛U�/��^��ޝw�<kmN{�!����òؑ�<X/.�����,'+�B�P6�佺ƈ�������sm�@~5LL�ި���/>�5�	����a�Z�Ltlg����"����k�5*�R!�����*oK)a��(��ߨ8��F�����7{;ڽ��s��I��m�֚�XݹO�uwv���~N(hμ>k��+5d�[�͋��,˫�����!Z�f�RK�����H��J�ӣqVvȗ|��ɦ���Y
���1��yʭ����hH_�>V[�<P7���a1��a�����.wIN�����'e�T�N1"�<�&�Gz�Zc�=��6��Rm�N~��,-}t�M�ҙSt|].�5������=�I�7�!��:;;nWD6b��n��gh�c��3����3�W��lCms{!r7�Y)Ũ��mZ��n�d:�������a���Y��>��풹�ϪvQ~zaG��^�!qe�[���O�uy?�2�� �?�8tx�E�+��xK� ;)q޻��GhgX�ͫ���0��~��f>�WT���s��	z/,���[�߳}�v]���X�̟�0p�ZW񁏦Mχ�Q��}�n�B���|��K�f@|��L^.�zά��Ҭs���*������yO����02��%�$R&F���
}*���F�q��2���lr/.T�;y ���:�Q͗�϶|��R��xRn?749_��+;�Rϒ��A=��1w���.����)4،���8��fC��r.�uи��$JX-"��oKY�mn���{�=��A�qͅn��"ԙ��l��*i��:��D�4������Q�5ߍi������n���h[�@��O��Δ}wĖm�`_m��f����V`h�������C�����w8�n|̽J���.6-����y?L�8�m�?3e�9g�H>u��|�H���R�~�{���4��18p��dC����V(,��-32�xZ���p����o�2���IB�I���庂�+�:�4�OPO�
�Ŕ&�>pV���*�L�FyZ-g�Vg���F4�"uTD��觳���ԥ^i��M1��<�d�,u$o�g����Gh�_ ��7ܭ���Y��8�0Ezܾ8o��)���b�W��}�k�j{�L����H��ݨ�{�Q�kˇąuII���
���[���Wδ�5B���G)V
���O�fs� �2��[���m�@<����u�DK.Y�����&j�s��=��d(.�/�yA��.��V�X�Ϙ����+j��]vv~UȜϫ�0�D�{����p�������
*�=,F
�'p�X�I7�9�A��^�R�P��y�f��vך��Tp�u:�Ή'=]s	�T�Uߢך~]1�F��5�Ԛ�tC��l��/�߄�+FL��~Մ&�3�3�IM�y�*��V<�[J�$Pa�Í2MW��j�����Q®=��R�	��1��_Y&";T*ag���Ψ�4����㠒�eq��?E�V
憝&�%�x���Jx�,��"gv>��-�=>��[M�zHw(�V�\8��q�ҽp� �i2�����.U��<i�%7� �y����=GM��3�.��MA6�F���H1u�b�z��W��a��r�FT��9s�w��z�X9�A��������j`f��M�؈��
SuY���l��!�܆V��wLl�2ڙ�c6ɓ�9�̹�6@��*�L���Βk�z�=��:���n\��a�<٭:*]�<�G�[0�*����S�R'�:�^�����2��㊾�����l5�/��N�y�X�.�0�v��x��=���V֣��zkL��=��ъ:�W����D�&�S,��4Do��Fz��n�r�	�ӡ^�ae�63��qyH+�~�$!��9��j2&|��-%�x�So��J���v��,���*��s�� ��T��w�)>Յ�9��#:��a�fS�j���:�S����7ɎH�ڡun{�����R��`��7<��d�R^u�����9����~��P��\NY���M<,��l �%4�#1�5���L�=��>,�T��+�[݆���<�{(&�^.=�+1����s�ݨ�*)���;ߚ��T���q�R��!c�rI���I�<ϟo߈-
��,��	��"v��j
!u���!��n&��<��/�W��>�څ�PK(yY?�p�v98K��s:��Tc0vI� �(�0�ô���o�P������m�+����/5�Ա�>c�^���������&������\o���d�|kQ^d.Z�X����}�u!�2�؀�,��܉�Z ��V��=�/R|��F��hc��R��d��Ѭ��Ng�!�Jj3��[�%vp�Q7\�A1��9�������W�K����f�uF%e�.*�$�����I�\*)Yeٔh.7K���(dGM�ΜK��)�\K;�â�0��ץ�e\��Y�xK�]���;�e���q����%�x4Vm F��n����/��$T�w/��1����r� ��"*��i�\*���#3��)�^8�J�F������G�_�l�:%��hE� ��&R
ȥ��~Z�P���f�Y��S�%גU*#ZW�9]T*�5m
c�����2����˖�Gvg�y+adL�e׏��T��2"��g�$J�~���1<�q���A1]Dep�j��"L�J����}�t&6�Z�<�}���H��.��~�n���#�;�eP�����+�u��#p�&����3�_���r�}�M1E���6"����c����Dy���YX��2�G�W����R�(/�?���0��j��Fwp��.�����n�������ƈ]�('��8޶%�h,��$�>�a1�c���E�_�-H�/T�,��Z�Zp7�.��nPW�BZȐ}��Sp��]g�h���1f�lCm���ѯ�<����Z���!��3JGz�Z.g�D6IX��o/��/��kf.���^�q�C���g�E�%u�g��);eNx�>�E�̠�������[��$8����!fĪ�l�u�zDt���VMqbYX(Z���Ä ?�%�r��}��CT
��Ɣ_Pv-O���|�i;5��პ��:ūJ������r_o��-;���.�؏�h_��xI�c ��ٚ�;_[�<��b��ݲ�"VyCz��5ake|~����p0{�O;��&�(/�g8��'����O����U麐�r�V^e71����w�jI6��Z������}U9���i�7�t�=���H��`�l�\�}ww�Z�I�'`�x�o'�٨�.q��#�;�q��#ŶO1�h�~yd�*m��Q?�6�5�i��u�:k���q��S�ѿt0'��A��i50_��J4�T�LݹshuWMpn����F�(�?����0����GC=sઃw�a����@�h{���k	/�tE��[V�P��Q����0��\e{����t^�e�Ѧ�p�R�\z\vo��� 1@p�n$���x\����e�˻��l Ā����A�i��D2J��]��#�} ��+ϥ�Vv��h-YSTI�h]���e;;����ߤ���.�9�ת����T��H����@�(�A���,= ������>�`:�5�9'/��J����y�sg�0w�586�g0�@�u3�'�t�����DO���Hk��kw7�� ���?YG���(�ue�P�Î5ߨS/��Q�1��e���]�-���%��`���j��Mc�f�s������.��*Z#��9�����֑ ��xvz]�i���)��[������h�S�+x�w���&}[�T��0�!дylurH)��"6/��A�U0��/�W���[�)�,��H {o�e���q� h'���1$AV����V	O��C�H� ��Σ����]@9V��g}�Y��x{鱭i�(��I�-���X�x��~�5-,��)�V�"���5�a�ZFj^�}�)Q��e@e�*�5׏�q^k"Rp{^[g���x� 3�ο&�������M�o�*��:��p��^�t����\lj�w黍۵����g��z����Gbp����H.Յ�l֥�K�4*g����yuQ%Q;H�y{�FA�K�T)��.�7�k�g�|[<�/+���;\	5�)"i��.Ԣ��L�p23��|�ǃ��콸S�����ގ�Rj�e����\ʦ���>��
S�|�&t-�^��aIbY�+_���	6fh��u�h�ˈi��~�\�E�5�V�.g(��)�������GcaO�^a�g��1�t�����F%��κCP�\O�?{��&o3Z(�w���e*�H��Au"�c�<�T<Z���%w+�3�?���MJ�6%��]���\�x�����i]-9�{�{z/�w-��S��؈p/�dM��/�h����uV���e�����@�[R����.��2m_V�������.=
B�oe�'�p�������(<��u����o��	�Lq�f}s�p�Cr�}`�f_�,V�$\�|��@����f6N�.�s�d�=�u��֠����s�N��ĵ1��Z���p��ý�6�X������TEu8��?�;X� ������U�7^����luU�B<@�lS��l�@p�k�/8�6S>�ٲˬ��u�{�{a�n{_�ڢ>��Z!v>ؓOqݾ^��K;>&�#z�	�J`~Ȣ�pVf�/�}f��f��$
����(�/47N}���,��=�nR[7}� P-�u|v~�����1Si�Y���=R�����͌3�g���5�U���8�����E���g�(��M� 0��+7�i���_^���s���]��᪼-�D!W��3����<*%b�����F#�,�Qp�P�'���eO�8.�����cjs�Km�eώ�/�=���4��ma�qN���Tkv�X�x?^ڟ�fe�(�!����*��FvrgCIġ�%�u����%�((���5V&_m��)�4+�SArx�����L�\��N�ѷ�d斍�b���y��<�[O��a�yU-�+COr��� 6<ݮ<@�tSLY9�+vĞ)]}�+@��"t�ӿ�rԣx*��2�\İ?��_ES�v?�e���Y������L˖.��IYi7N�G�B��\6���po��Wtg=ö��D!偖�T�A��o�t�$v����`� �O3���V�<rn<U���UJ�џ�?�}C�7��D	��ҨU2&�p�*ؕJW��2�*�g�ϕnO��
0��Ǝ�9�#�k�n�0���_m��p�OcG��<��	��3c;�)ߨ?��>j�����C�5�|��[��6|A���N�@.�D|ń��o<��V��X��/~�,%�p����b�j}n����F�N�e����i��B�xsX|ր�f�2�@�މ׼��H���-����Gx�۱�2�h�����t��ݲ,d���������ٍ��[����"����%a��`H8��]��ء#��@��Ȯ5��y�bF~�z|��f�ö�|��g���N��B��'?l[YU,�-k]���޲�{�>"=�i/�X��\y<���1��rt����tEF��tU����j��̫w��KC=�>#|W�Y�� �e�j��\JZ�O[ȕ�'�Tg���{q:M��975���B��8\^��-O{��wp@�|��Y���<��L�c�7��t�g��Զ?e��2���(�:'ѣ�?�Ԛ��ћ�v�y�ԛ�g���c��P������_��9pht@%R��~/��XK������aB=?��`�M̘��p��������1� �1L��$#��B��:T5��~\��G�F*�E���7���s �:/m���{�|dM�P��&��YhЎje�$y�&g��)���@8)�����bmQA�7j}�9�ǤZ,E�(�pkh��VHQ�Pk$���zJǕVn"�Uly�� L��gϴ�o{���43l�r�C*��4��4_���Pq�:%��PJI��7y�.�NucV/j�Q�g<�ft��MML$�i	�N�$���`��d��5��}�.���p�i}�-!Q��t a@sG�nSV��&�E��m���Ty�&�Z��ZWH�_r�����L��q@�U����b�6��6a��\HHT|aƪN�YƇ�8��'Ǆ
������mƲИ�_��2��Ekq\k��:���l������M��� �����Ч��!�Րύ���d����*��6���������o��|�>��S >�^��:�S�*2��{�ds#���"��7CL��ݒR��uS`b�xX�������c�)���e1N�!�9l|��g.SM�2����(��D)��>�O��`3�-Gl�=��K1Z͑?oDf?Q�I)�OL�c1��g��'[�< QAT��l�R�2`B������Y��0�˔#��m�� K�Ailb�{��}R�&!�b��vmPt�c���@	u0K��Ȝ/G٥��xK�:���!\Ut���x��Rn��ze�/8$��e�Oك�LsKl[��H����[2��G�x�Ҏ���aG��B;�&/���D�����W�wB,߮6>�5��r��!��~;�ۘ$]��������I�[J��"݅Gk�;¦\�K$��Sve�M��مuܙ��.p�e�A�a�m����8�QI���z��Zw�cI���M��Y6�;�����f�z�n`���筝�V��������o��.�TD �=�V�t�������;l�.>Ԡ�!��Xu�S���[�V�Yй$.V��G63�~�L�k5��ǭ�ȥ�����2���v	�/<��R&\k���	/_=K�gc~��H��/^(���G�׶�M�+_�ͰU��&��='f���.�HMK8aeC�-��t`9��r�t�c�c��������H�����2BEE��\ΘUq�H#���qEeBMyQ�Q�B^���u2�l�D*%f[���e�W�ė[����ބ��w�^ ������� �Qؽ\�yIOxY��W�@P �H�8�q�;�3��G�7���*=�5	@�l�Pg4����8ރ�d1e�IIM��zs=K�h��!0޻��P��x���4���+D=��=�G0c��4�r֭���3ml/����i���㯹n��n ~�1uݡS-OQe1MS/��Q���s1΀1�5�9���!� C�9V�Jh���G?G'��BR0;{�B�����Yp��n�c�%Bl���$��ᣤ���	< ��ܻ'�[�`�o} L$�hk|rHt�����=I-��\�~E�S��l�ߞ��@){vm�y�F�U�6��@�W��ɇ��պ��"	/ 8895�i&��S`HD��v������@��T�
�Ƴ�{�:��khi�1Ӽ��|����>\T��,�z�䮅)<�Q�@�@W���k���ܭ��z��n^�o��C`{*���xS,��軑��Z�a}�����P`V���µj�Jb�:V���	���;�(z
���`�[0~(�.��`�eQ}W^�X��kp=�'<��>i��_�rL�J���(�0�?���*^����\��b�`�/,�=����os��"<D�ތ癣ݭ����Z��Q��`�2�}mu5�a��P�X�	��RV��
i�ͪ6:|���8��1�Q2V��QW�'Mɼ��r�Z�OZ)=s�W��R��#h@�m:ѫ��j���<�� z�A/[����<����믅--�i�!��hvRRrb���K�M�.�T��� +�7��A���������q`-���)�n��*+�=r�m��꟪U1��i��hw���7�U���a;!1��'DO���E��*o�B�RT��������̏ �(����d�H�K.�ߖ��O.,��8ߎ��U�W2V933�	�	�-6���ϓ�)��(�kߔ/�n�ųHSgI{�ǉ�������˃//p��(^O�`m�t�ɿ�|��ΰ5���傔��3&G�_�E�\�G]<�}�=l3���>h�zF�����_�ȥG=�D=Ѽ�IF:��ຏ�i�UdJ%xz��W�����9�Dv���t��в'ɒ�����7�=��j�|T�op�D/�"���)q��-t�{Upѫ��;#��q�삑���RA�Hhr/|� ���`џ�7`�,�.���WJ���`�υR��;r������Q�����AXm�\�b0�S0������9��a���b^
%��."�:��	��r�C�	rD���ꝸ<����#�Ǯ��fGzerEOF�v(�$Œ��U��f_�q��sB�u�-�.O��/&?8:��E��BMIX��H'�e�|�]����Ħ�/H�S�٧��V�l�/��y5�sq��j�he��݌/��y��Iӕeo� ����1���gk[F���c���q�2��9��K�̅4N�ݭ�ƪ,�M�.�M��b5��/%A�y,��wGV�{,�GКD��-�&-M�.��n<��hv2��\|XX��Z�A����9-bxxx	<E\5� �ڲ�OD�^ť'��Ȧ���"p��x[�[���˲ӭz�C܃:�ٵHх��^�<���0+�56�E/�D��Ũ��8���*`0 ��̃i���ϰ���bb�+&�:�Y�U���LMMkڙ
E_��'�Ƿ�0���Ɣj��W#|����(�
N��A�=-�e�A��>>=�N>0>���H����v�V��	��0Z�$*�|��f�ZYY!N��w�	u�X�."|%�YZG5�F�hG>-T�Q��uwu��V�}�J���;���م߼�h����өY�9�*='?�V��%P(T�ULJ
<P�:11�[�_���?��0^��>�k��6RY��	���y��y��G�x������u$�7��kqU�p�ş0J�2<�^�nh�	;zӐ���=�n����.P��TǷoy���7!����d�k�]g�`��B��d���Z�qh��X^�� ��'�b1Ñ��a|$��lCԝԟ�OM�?;�\1_�b���j^7jd�N�y �-���x�A��M�d�zhϡ�9Ɵ��ADh�k�CZ�hj�v�Z��χ��q�=
,����������L�2˃XyM�8(G �eB�ج�o|��8謼���w�kz�����[7-�3�%�r�s�l�KP��_m6�ub>o7�
��#�Z�7hU��<�'D*R��]ID-����]��B�6%	�iw��}۲��� nn�&����f��D�������e�\j�ty��[�Φ)�ܪ�:�,�}��L�P����zY�c�ɥ.z�P�H�����x�#�������}=-44>��_FDn�6N��ʹ8Vv���� V8,��H��J.� ���|�g�5ӬH���mJ�WX�}��6̸�aFk��}�o��FE���H�B��Qsp�[��h[���e<骎!!�%��v���n�g�qjמ���/|� 'i�#��8��nG�`S[/]�E�$��']^��Lzw˥���z!ºa2W!;����~G��O=�����?}@��	Y�27\<�%¢Rv���e0�9��B�]��\����.ZLwE�c�D'��B�8F�}��{�F��g��Jey��Y����l��}GV��uq�'�G����PݕOW��:����G����R��T��=��kG�$�&&JZ{.v*${�{I��S�ӄ2'/�NWRSJ��;�A�g���ݨ-�����y�y���g���
%��R�@����U��z�f�9�����#j:����e㌲������9>i���7�z�=���_��p毒E������f�T��w���a�G5������CN��D=�����g����f���_��}yX���1!�95�3o���_�b'<MWfh'��-�y/�ԴC����af��s���R���>׫�x;�>(,�u7<P�д�1��[:!!�݉苎��/��۪��4mu��l�I���)�}xϤ�۸�.��d�Yt���td`#W���Q*k��X"�`�J������M�d*#uK>����rb�3&* ���)v(���fW�݆�����=WiIt��w18� �`OS�J(V����$�,11Q� �����&�fACv�|���p����l�~��Q��@C#����s64�Pr�������{l�s˔[ �����ZxΈ��L�ݦ�$��h������|g��ǒ��@:q�����n������}��#����=�UV�� ���Y󈉿J��8���$�����4�H�	�hD��v
�/�^;\ }X��N����\7�z�����<P��`���Y�
���iH�98��[O�ݾo;1��	\)Ml	��sp�[Òz�\�'Xt��#җ%S�b����6f�>��uu�tŦ�ݶ����mW{qo=�༴��2h�׷<��&�S�;:4eh	1�*ߪ﹌��\��lͺ��)z��0�w;�Vm$ ���Q3�p�ƥ��o�1����9�����K�c����Q�v��2%Ie�tl7���\���B7 ��a�?�!�a������ٖ�P��8����|�
���1=ey��#�%��O�p���)^f�+L�
��t��.�� ���
p].�L��f�{0�ż��@[�`���(DN%'>�;ʵ�?��.���LBЄ�����C|�t� ���H8���-l���x�B���s����>�)CS�O��#P�y䢧ݨɻ�'"��3��� $�|MHXrn��ˢw\��!Q�=2E��7%e�z�q�jr~�g��.���a�����Z����>���:D옟@_�n`OJO��z��	eD��A6�9�*C1�o���G��W��3�w������U�G�^���)f⤭�<�\xǦ�[��B��^pD����7�k�!b�/KA�_�^m��1y~x���KF�-�g��ٍ��������Є���I$Ȩ��P+�q��S��D�m���h�Ք�@ ��\��{0�Ii�Y)��sTx<�l�A��DS�g�}�o��~~hHy����/�(N�0��x�0�O{���9���@&s��i�H��I���)b#3�M�/�����w�}�D5�8k��z����u=%�u;��o}��%vrŢk��7/������_�y���Jּ�b���(.4���l�(��U���6�~��4�'�E�|}���d|��X�R7��lD�׊�nO�ybY���vBd'��mB�@ߔ"V�-sel�Zk*S[��h.IG���ąc�KT3ڴ�Q��jWrB4�c5*�N���o��I�D�>��״�?\����V���
�h�M�r�)�8����Ѣ��Ngۘ�$��$�PK�n?���C}��7@�^XL���
�=_�Zp��P�hA#N3��@<���9E{#C��I�"����v8���9�UD��<j�EeX��=����yl��L�~�z�7ڬ@���A����4�i7;�6VO?��7P=�� ��zB���5�m՘g�)M���|�l�շ��L 2������ax�V����>��>}J~�/��J"��#/"_[���@�� ~�rk��K���i���iưe:��?��X�`T)���Hm���s��; �k���!Oc(�����zb���+ybl�?��'4:tc(�s?��ٚ�|��cv���H�~������\�kg��Mڮ3	��>Ҿ�~��kKI�E��.�M��@Ko�e{�Jj2� �վ0�P�?Sd�+[FS�͡ՙu�a�!?���7(Ȓ8������K��x[^��o�o=u]?R�������V����U+�a��3�gJ��D�]5��GS3jF7�`lf���uH�Q���K*x�
C~]O�܅]�z��F�kp�ff�?�b�F��
� 7E|�7��1�@�	�C՚�q2vU�F���<�U�t���a��Ǆ��s����2ɀ����2��7��]�!�+o����S㍉� �''�<��k�_��U�%�`~��cgSŗG�0�/�u�t�3p��49m㊿"T�9����2�q��Κ�}��T���e�C��N�Qr6�nM��<w��eLp��z��
��I���{8��l}z ���3	�n�(�1@���3�u�[s�~I���􌱦�)�L�����@��ܴ�|�Y{��|}}�����5d3K�u�7�����/G1��5��@��_��5���^ღ�W��+C���Su�Zz;9n}y����:�W����8C��;�n�?�u����������d_G���Y��������w�k�w��V���wH�Y�Z�#g��;�*�L ߣ^����l�O�D4ey٩߉D�����В��%[��BsV�뚬 �q'��C�(��_����g�bʟO�q(�^okl��C>��4ט��x1l��^7u�vwݤ�C�;�Y����I���p/��4�@T1·]]��}6P��[�1�z�ű6}gT��Br���j=}�B���M�Ok>�_<���O���%%%)��LE��7�G����ݺ�ļV"�y�O����6wv���-�m��hXk-M�B�������ML��Jl��$v��<;F���Ӈ�,��bs��}�D6?*я�jI��Ե�RYI�/��� ���u���d��xe�X��e�;Q0������-�^	E���;���:���5��ıWYf�J]�M9V�\L�L%�������?Z^�O�_�q��ʗ
n�\V�������s��]W��.�ض�i���8�N�9m�>�������I ��Q(�x�y�s��t>���t����K��� S+x8x���u���o������X;E��1����h�Y�$�ϭ];��>�	@�C����EӺ�֙wh���.�]���T��B�V�H�i�����H��wO�ۗ� x� ���n���w�&�<y!��c��)Z��x�q �S�x�2��_u�-��iwX���27H��$ ���\q%�U�xۑV���8�t�%�10�E*Đ1����J�6G㵤gn���6��B����� >�=;�
�N�)�Fه[p��!�V��V�tL�{�kGW�/f��{rc+°�C'++Y�`� �8�����?�Fp�)�d��#,f����������8IKK�ى�

�f��9�+�G6���4`����Ht`
��d�Ϛ����E	JJ֚�����Tz�6�Ԓ:L�����{ ts����=[t��{�U11�D;��J-�C��t�!'�}n=G��)ˋt�㶑�8�:�S���^w�\;\{���V(z5�
=�@�\�#e� 47�C�Rb$� rc�7g����F�ͦt8fN��u_>�"��yQp�x��Ծ�mӖY"Yg$���n�\�<�'*Z������P"�`N�,��F穲��5��#ז�����D�kh��WoW��몖����o3pi���M�?^�W�08O C�ı�ݵ�q��췇�M^�;f���{���d���a]nݧv�^b��o��UF��BEGI)���b���4� ϰkS��ݲ߃G%*U�G�
��Tj5�t��zJ�ޔ���z�$~zL� v� 55j@�4�t75�^?�9ܲ�j�.��ދ���0e8�K8�p���%�;~N�p��Uw5���r��p�ȿ�|{��\JUT��5�K�Ąu��wBC�^g����fU���.R�i�_�N�^4��O������͗��k�l�Sq�V����i[�_�7z������z���w*���+MdG�gO_u�b%�<�꺱N��F�螣G�@P i+��@I�1%y�=H�������Z�7�2L�.��2��g���n�T=,t�-!f?)3�uY�t�R�9���ԝ۞��8 �a%@B]Nc����h
�g`���J;�Qnnl���/T�&��4�e|�;�+��2A�w|�q���i�Y-+-� hkر[z�:��I�9LU맔κuh�\�Y
��t�����V�E���>Mڟ�y*�^�/�h��׼�p�}�ۀ����ŵ������ͻ]��������R�?)(�����+2I���O- z�(���iMXZz}]�����~š���&4�H\0��CUM[�C[�����=�`�/i������������2�_��Z���7�7qڧBi�ox�O/1����>�uW����wo�il�}J�X�{y5X��M1��������~[��d��MIOQ�ǥ%�L�Ώ�ф|? \�"��qV`c��OVC	�sQ�ǗkQ�;q �Ŏ1_�[�:�GNn��ϟ�3����$ Q�s�?`E%�)൮#��MRw>K�Ի�K����5U�!�OK�J#�Ȫ+�a��Q��#� �w��m��+���/oX*��2
��O�.}
qt��L���\�E���X`�o�i��������QQ�_��H���� �݈ H7H�tw�4�-=H��R�]24Hw�=�����X��5Xp���|���{i�;���c�.��n���,Ro�J�fk-��J�m_G�8P:�+�k��0
��z�D���cn	�z[q`ٽ��tH�����ڔ��/t�{0�,�=�Ck ��n�H>������:��ѻ��w��7ʪ��'����h���e7�tyqO�C׼p]�v2��R�y����������511����$�ˈ�i���ƻw���,�|��,<=S�I�|�������N���3Hm��6���}i� ������G�W=$\2$x�#��J`{��N:ۃgX�>��HY�׀ԟh��WYë�hP���j�!��<�m}ML�e��gy���*�z�]�;O�M�!Ȫ���Ի�yf�l�	���,��9]s��ۓ�X�-�Ow�jV����}�y�U��D0Qe���8n܊L�\~C���?� v������6"�	pa���������?�3���X8�O$R!E���V%M��;3�7�_�k%�p�.�﫯�K�'ةUe���~��q���b�z7X�J�VU9~>��x<�\��\�L�ч
��h�ri@����a������pY������ZU�0��sK�A�=�����Ő�H T��! ����� *�-����OOmmЯ�ƺ�Sv����V��|�����uR�k���m�4�b�!9EDY���J�(�z���S3@1�lK��E9.�����];[69�����p��Bm�����r���Ђ~f��;%\��Es�OF�A�����b�,SL�i=�i���eqs_���(��g���(���Fb��3�=X��O�LYC!���lOP��Z��83��l�2�8Q:i4���2����<a��VO���.����&+���"s�N\
UG�S��݋wR�m����㬭jj�y����+���\�*�Se]��A/H�r������ĺG�B	d�A8��c21YGxn����P��Sl#�px��5�/8�ٔk;TH����������]��:��Ǜ¤�16ğ��4��W���E��vaT���B���j��H�>����=|��jjv���#I��Q+�n\�j�TWm�4J�+���?U1lL�d��.? ��j���	��o1%0^e�u�����o�>��b�H.�ߓ��=�6N�� � �Ι�ݯY��Ϯ��q�ekN3*��a1_��KMÃ��LS���*��dBv��p�n'������5��`�2_����B�[��y�ns���v���ߢV���e�D���~�����&����d����>y���q�� 1�g��ƸV��tQV���:����n�Z$s�s�k.gb�^�[�h�5���f�n��o�W�)�:D�T�o��l{��n\�z�&�眪��Sĺϱ��3���s3w��㚿�%4g��]�=X����|�t�j��5��`�PQ�͉�Ԃ��Z�¡�b'+NΟ[��uC��'r�c*l�		��M����
)�����J����US�	�dZs�c��^<��c~gyh:K�J52��dԐ�д�����V�pv	$bpP��� ��pƗ2l\Q�����+�L3 ~RǏ��h��t4��Ŧ]O�lQAC�,�16U����K"�?�ų�yb�۾�n����YD�6Ɖ���;���A<�_4�J�2����O�]���-X���c��R�Z��/R�Az��lߌ3��������4B<��3�;}��4R���T�ux��5�"�'*#^O�g�7B��׆�/z�>�������@4�p�@~�8l�L�)2�q�DE�Ţ��'ϡW��U�|F�UQ�oP���ob�S���c]���ը��m�X\��Ax���'�?*��f{>�\��;�t��Yƾ�����$����!��]1P��3l�Bz�&$$?�ۙ�}U�$Ϝ�r�r_Ub�C6�'"eS��T�T�id+���w//���_zm������/��Z���v�j/��Ч�C�(5�5��yƦ��UoN�5Ky�]5n.N�mOw	�������6Aq���s����
�mE��5��G�>e\���Y	Fe	�w�%��`�����7��iD�|�\���>����*�A
��-���G��O��B ��@W���9�o�'t<;�E�:I���q^�4�.����w�1bQ��9
� SX��{�/�F�s�"�&��������qr]�+Wttt;oN�N�ZX�8e��C�ɨ+F�w�f�0�qk�Ӳ�1f��^��e�% ���WK����o����F���	� �9QҩS��9�;o!ӿh'\<�$j���ג�:;��5�>��_��s?���̆#���ߠ����G����"Shf0�ve�^���S�Y+�*4s=�0{B��dD��_�(�T4�PĐ�YurJJ�����BLL�
n���
&h��.F���rIF�jt��=�C�ʾ4��:����Ҥ���C��ސ��;'�c�p��]��R"RR߾�!�j��	���Y푩u�X�G{����{�,J���hk���.���������8��֖o��\��
��+������QZrϣm�^<?l'�0��Q���n%s��!"W�"��M����Gc��Y���{WBֽ�&
0�J��ތH�2\��`�X��n�[ėR"��|Q �P�H(��7ˢ2D^T�\W3��/�}����-)r5��2>~	s[�Xӿ31����p����z��>(����6����v-5�tA�V��G��("a�G���t�G�K	g��%$��E��=K@��{���TTt�+��!�VFg��1>;�.N
E�T
�K7�=��q&b
�l�u�"��}��>#{�<Z57!����н���t�Jw��ۖ������U�'n�il�ET�� �������Ky��~^�����ϒd>x"w�1�n�z;s�� V��"��"�5�J��i(�q�ˁE���/�Q���K�_��K*(`�2�44�#{��w�����u��S��_�vz��ccc2w��b��a���"��I����/&=��'�5�]���:���
VJ�o�"�Wn.�/:Dn:L��+?kNp9"gH	;�!��)+�)�2��w}�I~fS�թ�A�����s~�ޙ���J��#����FB�OE�����9�_8K�^�9�޳���\z��sً�&X��ћ`	@"��������Y��#��
���[9q��&�u�Rd�_'M��c�;��4ajj
{|��ѡ�h�Kc�ڀ<Gv�.�Z�>v!��B���|xl�ӑ�l�".���	�t�%S�;eJ���ĜI���NQ��K�+�ٮ�z'ۤ���o��)�}�/:c�U��ĄC����uCƻXt��"�y=�w_ J����v}���~����Z/�AdNgˑ�[K[,'ҏ�w��~���\�� ��C�6�7����^���M��ԡ���iHL�b,�\I����K̟�q�"ݮ�7��=�b�v�D�0 �GҎ.��V\_�{�͘U���R� >?���$Q<�<�G�7��8l����ˋ��\�>��Ҏ�+��y��)<�H
�:\}��F*ɹ���uJ3F��9v���F�֪~~��s��g����C�:\���>JK)4����q0<:�n�eʀ���L�#��j�A��E�B��L�mR1�a�S�wT��{����ɚ��Z}�z�@��c�X�pJ�V��ML���r�VDU�.)i�h������^�������׭O����B���\��1"��R$N�J_���ȊEGw�_M	�u�ϛGh��.��E�b"ަ�;�y*���"]��!��ၛ����ʈ�O������;���6i����OTp���@��5��y���N��?ے��k�	�)N;;y��D�,�5z;��^U��N��_�M�Et����q��i��|��e?5LEN�c.��_fF�5
i�0e,��)��BTD$C]�a�l:x�ͧ
3�X.k�#��	,���D�c�첅'������"�Ps��{�}�ފ�nӋ	#A�5�Q�m⓬�3�D�i��J� �!�G�w����6��x����|��^9�h�~.�=�������KӏÛ���2����Dz��w�r����Gk�G� �����0&���+�0��.�l���I��s�FNV1����`U��h�����p��M�B����@���V΋���f|f�o���?Ǆ.γ�n��2�y��OuU�ڳ}&ː3d�E`	}^��ó�}r�>N'�7؍���x��]�l�}@��7��I�lez��i�f:\ѯNk|8�O&%]�PL%�$��Nj���®F��
�w��.�~ɉ6+�����\1f�c��]��\+�˰`����l�̢7c(A�4^��n�i�~=�01I:5Xe�$�ڦR��~�C��݊%n�d$�ٸ$c����U�.����o���Om�0y��~�Y[�ȋp�4B��a?��Y�?�z��~�n��?�}���弯/�60F�sI�O���E���/~��o�{	��`ϻ���^�ę5�@����	Cb���CE�]?>E=d��c\P�hr^��������/�b6,W+0_
_��{��'�<�e����U�?�mʦc�/��9�p���uzk�˥�2�«�����*���"�qY���Ƚ(�+g{��6�ܿW�9>"�5��+d���~zU�'�#4TȆ�\$|<��G�M��|g�P�����2��czD~���1�W�(���]�����3�J`m���2D�����S�scp�D��2�& ڡ���k��������
�E.zx����s�5s�f����v-'���W�c�g�-���v��a�A
ގ�w���kA�
5��Dl��7W��w筧'��7w��V��=>����{��#n0-z���[|x��𘅸��\���c��ӋlE��-|9,!��G�
�X��+Gهm��\)9�>��@��z��Z�6��H}U�o��_DtR2�9�^*Ȯ�g�Ǽ�@a�\��z���#�c:����A��N��� W��h�)�����r�h�RS+_��U�Uj��:2j�d�/��4��a3����:l>q����
xB�G׏/�c �_�ίs,&�VX1���f�	Rd����5���;ׄ�q*/G����Z���h�B�l6, ��'�5�H|D�U���R{����5Ƞ�����u6�qC�Ƽ�窢���������+�q4g����(�Vjb���5��ev����?4�:A:G���悼	�����w.���棍T�~���q��1~\"2R �/�~�5�Ԝ0lz�y��G� m��K�i� w�K��^.�AJx��#Q��]��'��%�+צ1?CbE4wx}+�&>��HQ�-��o�89#�sgǺ3WD�#B���U/�SY*B��-�*���!B�}�:ZC��%*�W)*��z����䴴^m9c鋝���:����A|�n\8]�7��qZٳ��_؋̏h�T�%& �E�rp7�(�"X�1>�*�Z$��R���#YɨB�ƥ�)��c+�tZ����_5^;����f6k�����܌��H��>�^�::k������'ZkST̖�	t���<�hqb8@WW5�d!K���lH� �7-��r���'T��z�����r+9M0~)�
:h�>[�G������{�J���TIWW������2\$-����B˯�ηߞ�/�6�%��󅉡�ll.��p��׏s�˱���.'���m����#��'��A�HY,���.�]�P��Ȟ�0)nlF��ٓZ|7�l���#h�t��uk^��aP���)\z��XO��,����yv��׫~�Z�h�H�����v]�F\>�嶛�b>^�zj�����A_"3��"��`|lj�'��@\�x'mK
��a�o����Tgg2+�@6������1��łW��5w�XЋ�X�Mܤ.xT`��l:r�utE���v[+���[�{c�uo���������KՌ�׏U�ʦ(RR-���X���d��_C�'ss����>�,׷D��bff4�_��"���l�oT��eoi5�����&�]�����6F�&��C8��(�D�S~r$	���������]�A/��X����G�zu����D�2R��J�c��kw5iԀ��h�j5��W�o0}�ND�ד���U�������W�̇i2Bw"w]�PH��B`c�MU7Y��4� E2TI##���+�7VO���X�:u�)h=����鮪������2�/5}c��*;�X5��ev��as��/-P�ְ��5�����;侓i[$c\�urv�\�פ����2޻��As��{���9	� 0r;���:���D����iY?~�w Ʀ�N�¢�u�<�j�H�'�lCՖ�����g��|��ࠧ�?4	%VVV{9�����L&%r�e�8��H#�v��R�-�S���g��d38��ߖ��8qCmS
�ݥܔi�1{xYY�g�dM�����s�J������(�Q�����z=V
�"�ok}�[!��_C������t|y���3��N�b��"�adg*��.֦���궻�'D鑹�=e��D8�^��状������_S�;��e	�wգ�H�}Yi��@�6�<�������*�./��6 ^־�Pe�Ƙ����At�S?� ��7���*�!�y5=[�F�\T_?l�a�QJ��
#6�����pu]t�/��)��(�1hZ*�sg�˩@SM���S�yjH@ \: V�INcg��_ޯ}�%~.'��x���v1�_�f���.|�פ]�lw�.��>�����?�H�W=�����X���~%�Y��W�gb6e+'J��P]天{)۾������#\3]h?b���K/�X�5�l������Lu#:�H�:��W��ل��m�����Ϣ��k���﷪Dx8g7�O��x�
7'�3�:W��`JD�dݕ�(0f�F�f�����hc7��G"9ش�JW���?��#���?3Q��ظt|	��{���a��#��H� QfF:�w6���o��6Z�rE�*P|�o� 3iLn>ЖF1���%1@tF_�RƓ��?й������'9qY�@�(<��:�����=��9�غQν�ڛ��5Zy� ^�`���_�b��v-�������W�j�ou�2�q��hf�s(����p��ʫ����}��h֧�f�zkgǂ'���I,�vv��w���x۝��Ү_ ���Ct���`�/>|�^��	�Wo߾@e)S$|�U��|��Ƴ�gE �[��5�/7f�;5����&!!�k7v��d���":#@�2B@�P��i��!�]WJoػ���9�%'Һ}��42��k�4;Q�6AJ�H��򾖩]6�RT/�]Hj�BAIU	�r�A�@�N��(Sd������P�]]�k2~�3���_��L-x����`5��q~���h���F����b��<���gg��aj}��"�B�M�ڂכm�2	Ȍ� �"O�m�M0�	�R>G5�.��z�w�L0<)=�䯨!�}����Ԍ��Ы��E������81�8��p�t� ���Zy�x0��w�8�Ԙ�qqh�g��M��]�K?�ڔ��V���5����|����{MM�Yfy�sx R}pN��Ki�|�ϖy�[�qjjj�?F� ��I�õ��6�G��]}{�)�?�����ʿ�"D�Z^����[�e`��l(#:j��1�ȼ��ڭ�+M#�/�ܹ���坑<����%�u���s��MHϐk���^ �K����禷4"kR"ᚅ~PG5�|q�ٵ:��h؁Kn�x`��׍&Y�9�L�'g_CH�:5L�4��2�e�xz�\�1��TX_�	wN�Ӎ���ߌ�E�t$�;��@ԡ�r-/��^�ϸ���z�8Y����T��5����{��e��ܭ ��F;;�-dK�V�̚�(��-�A�Vu?�
[a5c��fh�0��Fq��(���0�y/�_b�8%���~c)��E�]_q���g�}i/�l�y�$��� �ky�7�5�:j��k�!��"�H�הo]7˃)Ajc�'2%�Ǔ�3������+�1DE�|6���㚅&4Y;2�'�!�$�Z��0~r]�]�kDRΤ
��v�t��G�z"��<;9Ǧ��=2@���Ҵ���jE�KPH��6�K�uTw��D��%F[gR���%5���fa��~`G�=��r�����="Y<dھ��kV��Q�{�4}�r��"ML�����ҏ��pF_=�.0#��5Z]|E�� %?�c�1�����=�6T���]E]1��M�`h�)��t����;l��ݳ�4k�����0;&�w���Q�d����7-�[zܜs�3�1��MO$��<L�r1c��T�\u}�@����,��U{bgܹz(�\a����a"Z�s]����dh�b��[q`���X��W8�u���Ӈ~��Xx��Ժ��A�%t	��(�9�\��8��ޔ`�Z�D�a X���w+��""��G O/�JTJz�J��p_7HЋyבb���(���c���۽�cX?�Ci�ٳ��A�}7�oL���C�}﮲���',B���-�,���������'
.��a�J�[�-4�d����aA$54Ԩ�\�B�8He��tb����kr��U�;x�K�y4�}��e�Z�xy9l��!?$�t�$�$=Z��d��_۱j�c.n��0l�{B�����PR����B8����-w��C�c�w�?|�6It�\�n���#���:���|��(�3�b�Ю��wY[rսYUWR[��A�vu'�_M5-�|�;�gh�?�����yuf7Đ<!��0_�Ȟ[t�g�w�q�vrZ��#��!Q��m�YO~����ֱU��5{&��!������+�(#xA�Mw���8Q��`#�{8۔7�:�HR������Uｆ~�!�߸��w�e~����	�T{8ʗ�/�ł�x3�Vt�Nmi���ô���$$�(��/ϰ~Rǅ���/l%�F�|�T��tk��\�D_𘛳���c1��Z^hh��e�;/��H��j�����܏�֕�s��wW���w�[o2�K�ھ��tҎ�L�9�ϖi秋��{�����K-n��y�L���d�8��[���v������9��þ��!�c��*zI�Ym�nw�J�tuZ�?Er��~g�2�L���>�`��{����1[��0d�n�ϗ�W_y�Z��SE!�o���v�yTz$�?M�N�hV�$���U����8�-�������y�}�Dj�Rh�.����%���N}3�c~'�wr�8��2mY����������濲��O�J����^�6�*�>품�=��(����z���L� I��	���`dܣ��f��w�*���,�.o!6�(� w���;�f�r>>~�w����Ǜ�u:�P������pwe/�����_�䛱,�,��5��j��ɺ��x�pa_����T�$�1w���]���e�tr��U(��3vJ�&-Gę��� W��}�sњEV�5�p�i^��5��hnqm��l�K���ϧa3��{�lpim��l��LA	�H���v��jԿ^�DL�Ǝ�̰�b,е$��j8-��T݂�g����@J�%]����qMJ��;�/�{�2���H@�������C\�m�{�?\�G��P�B�}�_e��w8.�e�7~��`b@�4���o���P�}�i���XѬ�^w�}�j��L+��o^�\�
�G�s���(��H��퀐l>(L���Uw24������b��tĽ��K�_taPy���جLe	���b_s��?�a�߱'޿?��K�oЍx=��Kv�Ɓ��4��P�L﾿"�a�$�1X��^��M��Q^u�bVFS��t��n��1�[�vU��Κ�{,��=��yq������Ⴂ�|��	�5k�I���&3�4��~>��|]B`�l���8zS��j�����R,�Q �5�̧�B`����am2$q7��:cA�|�:&�g�9���F��6�KIoy���il�EI3�$�G�N�_�y_�������l�d��!�8��*C&���Ve͑v��U`15���Vc=��o'kQ]�zL�֢����<�	3p.�&t����Q�9�S����@r��P��{���w.JΡev� ������d͜��M��|O�v��x�&�h��ͮ.���	��֬Wɿ4�~8#��Hڌhu�}Y[�BҼ� rV�����u�K�.Q�7����Y��`\��I*��b?(?wJ�~J;�~�Xٸ���j�����O�3ow/o]I�7�Ԃ���Q�&S�O'`�
.Z����]�.鋴\���ؗ���`���n-��7un�H�XP?D��-P����v�ц0�)C|]Wdaq�o��p�S���j�;�� �}O������ɸ� {�njY��o�;Q��'�F)�_�Q����B�3�NK�6��G�wϦ����L���������q�E����l�i3�j�ژC�����c����l�瑟�C#迃@�����׳���-�m	%�0��1�~5Ta�Zñ��-�<��;��L�V1y�i U���e�g�"e`�8�o0g��Kbq+jl.��Y����7���pE��;���1��*�.��I�A��%�IZE�ngc�s����Ǥ?�D�ۜ�f7���5�4��S׬-!���t|���̀ϩ�yĹ��5[?���8G���Iş��]xyh�zY�cu}D�Jz��>b�Рv�'\UB#�q��8�`���Z��9ҟ<�׈��u�����-7r+�j����yoq^��l���Y��ۙ����E��SpH�%��+|ks6��� �8��X�4���W��s>��*�����.��n�O��8�ķf���H�[!�϶��NT�d���$�_��ƈ�T�}<쥅h���3�?�5�F��S���fw�� Kg١.s>�g'�si޳�La��7}Θ��� ��y����|�_LOG�x�{�9<JMVa�{$��jⷧd�igxyM�FŎwc�
i�߮�@�ީp��u��Ǆ��Fn
('_�a�9F�������P{��@���'l�YU}L�.��a�]�M�-��K��.�����I�-j���0Q@Gv��ז\r��䞞��p�h[�_�J{;��e����=%����l��Y^9�+	������O<p�s���h6�"�{u�����1�'�ô�G����}]����A�����?>5b���n�[t�~ϊ�������
���dcu����I�e�Ϩ�,n{��U=�'�I���F�E�ȿV��%v^�� �X��օ.�~8CH���|�������ˀ� d^V}� ���כ[#փ]
,)��:ߣ��6�aH��r�_&�����a�2���4�Kc���Hz9eJ>�}4�c�"���0Y*�7���{�n�MXq�9=�-@�VZQR���h�/�{�8D��0�,�uw�P�����Ѥ�)q):�|���ð���	Gyj蓇h��4y2��b𵮐h���I�B�������"�x/ݓa�������Z�k@��Z�G��	�3��k]��0�?�6no��3��l�2�hL=Tk�A]xMf��O�|>��u�Z�%�==\����L �۳H��y�e\u����V+��ǝWBf���^Iu�_�ʃS���J�qQ&�*.�E䁶W�tp
�I_�4yx긃��C������,ѩ�N����5M��9Q������������-��
�@���l���Fr�C_���>5jRR�����XU����阬k�{�ǶR�˓�ۗ��9}�R\���#��,_wʙR�`���;Ƿ�����0u�	�Kcxbx��¹��1����Z���wv���@�[����ġ����O>�T��\�K�=��av���S.�n��%e��P��W���,��S�s�f�B�Tm���N�޾j
Yh�!jk����y$;�o@;;��N{!���
\�u��Uڢ�9o1�T/������ZZ����V�ˁYtX����h&l���@<I7\)$�xʢ�^�vW���=�3����O�a`�w���H(6�����FK8 �C��������'��=���\�OhJ�4�FEq)ԝ/��޾柭\@�gSu�̘��'n,���٤h��W���,6����;�/dFA ���#�\k�혣D��.��U��Cc�5�ARW��Y�=��O�������/������-o���A���H��QNt��^��
��<V�*��a$ �K��ۺ=�X縷��>���v�����o���$	4�pQ�sc�[��qw���ߌ��-�Kj�.���˧�̩Ӛ��B~�2/P��ʗg��!����!}�Ãl�w�j���'�K�=)囜C<���WFng�`.��˃����%��u�ձ?�_�����F���ξX���̝��G������k�K\�lK<Ǫ��r"�A���;��=�S=�.�M���c+0�n���Ka�AvS�G��m�TI����.@�C���䖦�f��k;O���k0'/*��'�K�0������;?�y�qlk�)���k�Mߧ�"��F�9��<jD34n��H�ˀ�*��Q"Z��t+�W�%��63���pѹ����H�K�VM�<C�t�o��Z�墺�
ɧ,�IZ�yET͚P�z ���O�E1/����7$�GVvT�n��F�&�L����@��j����ۢw�&)��pA������SQ1Q���j'EF�g�����o-�����EQ,V��"��vm'ME�F'���{=��w�o�~SZ���x>�+sn���3ܻPB�o,զ�/j�m�d!�t�m�j ����B"�R�<�.y�����>��V���~���̛��8ʬ�U/�AI��?i��x��o��5w�U� C��⻝C���o�qpWRNc:���v�ը>�`�XD�jh��W�V_��NH��b�1�Љd���&�&7D��+�Hݣ�� :Nc�����3&>�e [L��'���@	����K�R2�)�\���g^>U��U���Yr�|���|��ٚ1G�]C�n�D�'��F�@�� �i!�wX���i���)����r 9�F+�#T�h6X�P=��1;��uq>�9#�j�!��kud����;L8�s�&�! ����%�"�Y�B�2	��;��_�fVlu�tŷ�Ǫod�VTl6)��i,�l
Ig�6����k��@���;O�� i��V��-Z����Ih��vd� ��E ��X���-�<C���� !��n���2�߁vf��G���c[�$�3��n����Y�#�����E\{����A�ƴ�������)6��Y�%F���!P�5�K/�p9���l��IG����dc� >�����-��^��~{������r�}�N%��٣���k������w]��('f!%�;z�fCi��N�b�i�_��
�7�k��|/��W�Qn�6�W��;���&8�\�3,�%m��{�˼+D�奷���\����C74m��;���r�[,c-~���.�֓j���F ��t3��gng��-�cZ�uק@��cHjܢ���'}]����I��lV�����e�zNp*i��6�,�S�+*ixMn�!m���I��.��(���^��+��:�ax�[��wx~�_UOz��'�L��/���{@9l��X�<F�����h���/糛��;U<_ۉ���r��� ���5�V���K���3�H��ⲱ0�լ�P��m���{��!������Qjq�$�`�pM�J��/)V�p��2�wH'�����Zal�eA��)=�R1�}K%`�C����6�?�S����ߠ�~�Gb�J��t�c!����$V���n��L<�yxl��)�\���i�U��E[��ʚЪ�d���i���ހ5���N�K�c-�?:� ��KRW�pPU�)v~O@��������M�R<�Lk��t݉�F��nBLA�l��볽��]ܔ-�Np�Y������]Q�Rwᔟ���4M�3е��4a�B��u��Bny�-����/�\�byT�*����	�	�]�tC\Ѩ��a&��;�͸x	��%���w5�������5��W�8p.v���U��[/]旷�N�)������R�u�����t�ұ,o���KX�ͨ�S(�\"��c�n�㯩���ԡXr�tS����eޗ�Β�J��C`_-���%�}f�iRM烤��.{(�J5��	�d#�
�@�ݤʭ��N��Z�A�X	"��cMb�H��dcĽIdt���c���x��Й�|�L�n� �2���WJ�6�~m�#m��p;{c�ǧ��]�{I��y,)�=<� ��-22�i�(��ä=��ܰY����om��@q��ޞ�T]t+#K��v�[��]~�Ud���`�k.�����T�x]��hS��:{9�nA�K+�R>	�eEl�Nu��V�<R�0|"K��q��U?�\�Q5���zb��,��0a�ݭ��5z�#
!I6�����;��{L�k�a�Q25{��e�wH,R�H�D�h�[|	���=%L��jm�����A�'��ҕN}��"�V��a�>2 ��Ҫ��CB��z=�� j���ya�&kR�/ooKm�t0� @�7zDl��l��B�wHF�\L��O��l�Ko1�P�~}HN��}�"�.(Y��W�x5D`���EU��%o�F��f޴  ���y9�#7˫��d�:��g��t��(iZ�`fH^�X�������]K7=Y\��IE]�[��@�Q�@��ŝ&RYJ�6�\�I��X�/jjN�$W��ݺ�/¯17���d;x��D��@���9�t�����A����moF�7�7��b+I�߾^�Z��	hw�=�M�o�B���`�?��茶���h�rH�\p�[�o����ܼU���|�xQIͶ��_EM4t3�7��C3Dr�v�s�����<��n���I��� E�sU�\���3�@x�#�[�b=�-@�2W��-M@@����������})��^����d�ffeZ<��5[g��A�/חlO��<��_<�g�t�̹8�������䊨��\���H#{0)O��
��\lݖn���s�!�\�A���7��)�vj�C��^��\��Ms�f�lr����,��:�H�7a�o{��F �Q#ܟe�aͯ�"��]�?�|�z�>H��=�F�«��O���jR)��GH�����{D�/��Y��J�(���B	��"����^�&|u�Ҫ�	�] ��bi�q;*��|Q���|$�PD[G�E�Ւ��*�z�����͸06�E���q����l�uƎb-Vj��i̬��XX��V<17[�L��mh���9N���uj��5g�Q�J���q���@z�k�
65n4K6M�eҍ%���	G��E�򾫠:`����R9$�'�~u���_�>�>u��ܲ!9�ȩ6ьr�>�&��ۗw������[��\J�ŋ;�w4X�{��}��Y�U6'�L��CP5�#�=�3��$�0�>�O��/�ْN/�=�/I6�9��*��թ0"�kjsY��+��KY�C�AB�❴�73��wܳ���3b~�Q-H��
s<��C�����`�j�u��ؠ��V�^���
�$3�>0�l�/���y���&;��J�֨$CS˪;�� ��]~�d�2��	F0-�Ju����qjrF*�N���qu�]˔Y��)����b��
.��i�r�0���������&��9i_	�Ƀ�J$;9�w ���:�8�Ϝ�үo�u%
4���� @�.�_��+���-[ �6�P�9�,w�I$�C�ԉ�n�)`�"P��r?U�����%����Z��\�ڑ��Q7����<���q��n�hn�}��sF	��mئ��r��] r�xm����NF/�Z���,�ԗV�z�.�K��D_�^����}�T�=�4��er� ������ B�83��B���L�"�0����v�jW1c:�����II�������x�M���FQ��W�����ȱaK��'OE�l8햿N��v�&ŋ���{X�g �����^֨F��F>;����?���}�hK�����آ�yh,��#P�O�����"x��_�[-����(Z���F�t�x�c���He
E�͕�b8��u�ɭ�����*�YW�o�S�y.����N�ʸ9&�ˑP,�H�N�y�>Q��+�����}c��W D�|z��h��!jӨ�����	�-f]�B�X����V�l��]q3���U���^�޺�ٚ�km�f��l��Q'K����=�����Ugꍽqo���$I�e�W�\U�ݐmc�����7�<� ג�2�!x-���_6ate�$uHj�]?ۧ�í�A�A�Z�*��T ���:2@��N�B���,a*
�����a�U��]w�ԯ�iS[�p	���N�:��x)�Ukw��U!`�
��椭�7I87������<��p&!(ե�G���|#M�Э\A����G������z��/i�	��|& �
��/����p"к��^�'į�,Z^�kv�Q��y^uT�����WV�S;���3|w���
֨T��o�Qq�0���`8�_�0hW�����;w�u8f��R��־�����\�ͻ�B�r�e�1�qjer��� q�<�?���x��/>R�[xK��BZ��u,QYb�,Y+��o�0�T^	!d;ٓe��P^�}�i��$�c�0��jy��<���s�s���=�޹���d2uD�y��P�[fVU �/a�rh5#�L4�zE��#0�V�p��L�az���К��!_h���U"������3|��#���
��<��s�_��:��2�n��rʳK��3�Z�C�Ip���Ӓ!rZ�ּ�st��UՄ�w�ӝH�P�;&7���[����%�U�s�~<p�Y�aq
O
]���-��	�<�_�[��m��ßj�V
Q?��q��3>���,9�iL�I��~˸��b����^�Ѵ�����n��/wiZ�{�+<��Xf���j]:�x)�����p��|�Q�q��(��a���:r��i���#vh-0���Ǡ<�:V,�ʀ�#0_7&�����*�q�]�F��r�h�&�����T�����]�u�1�<���2��7�>�{�Ԣ�c&���	w��4�J����G
u&.��M��G����ڎ�6�صZ�EN5�Ϭ�%����)���տ׻��䶴$~�l�޾��m�ꋰ�-�Q*g�<�LX��>�<��m�y��޸���e��]k~~��28��@�m�X%gZ��lp2�x�^s�G��(�ҹ��@�`^
?�?l'�#t7�o��;
~s,c��F�ZWՎ�����3��fX�D�0���������2�fB"���|�5�M���F�����;�0���5u����jaч�����@�4�[r}��a��q��Uy.�R�vˤ�F��N�Bo1wϡ��3}ˌ��}}�ã�;����hR�HE�%��ʔEig&���0�[QͿ�;�W���؉WW�S篇���[yQ�a���}�t[�sY4n�NUU�������L�_/�o�Z�m�.�p�����Ғ�ө�1�,��"���%=w�������t�e�m��V�_�܁gV�)Y�nח���������q$<g'!Ɖ��l(�>U��i��Dm�ٲg*5i6��XLM���E~"�_�E�e��TMl���s5��I<�B�w+��c���<u����V�3�:���Ū������
o{ԕR,��q��-���3��}��8�ޮ�yʪ}��nHt�\�.������#�^�W%��-�n=9 8,&�M����YP���q{`>.�g�8�S��w�ߙ�q��2��򓿰Ar�:���fN�"a�L�Ӄ=#ˋ��D	�c
� "��A?-w���}!#�&#�m)�r�j�[\�)Ύ`�!�2���h;��;M"��-�K��}Y( �H�&���7Bύ��S�V�<'*Y�M�sJ0��F��~G/����^|ǧ���3�FE��ִG��V;k�3�i������C��+#�O�g��y�-��$��
�R������4��v�Nj�{@_ψ�uR��Q)J���>߇���r���K��k��b"Y��Wޟ]�, �j�^�F
�姖�z����殸ڄ���M.��j�`{LC�@L�N�D9>��M�j�M{pK6a'��m7�9�!���E�g5�*��.ÿ́dW����Ry�P��S����_����K�'0������}���<R�"�R�ղ�\�~(�@�c�ϐ�[�Z�Y0��X��`&nmWt�7�)Dy��Qz�0R�q=����:���EL�Q�С�Ɏ
�ӕ�j�*��{��y�ܼ\�e)ߴ���W�U���j5���3������`��\]'G_�G(S��BN�����_�PQl�,;��)���Nr��n�6����:mf�}�Q"+`ݪ����M)���(�nӃ��A9D�Y�%[Mx���鉿 �o4�z��x�1}ϕ���d�:K������v}󋚛�%�%��i�b��;��rЉ=xp���½S �����$�W�0��K�)�(��q�������{�47�V��_��UYc�^��Q��}���G\���e1�c��0�&fͤ�X�s��ۀ�j3��-7�"�(:U���S��U�8~�O}�_������2�mKd�<�D��T�mu�*������ot� _كoA��'��A�ӢsE��!�S���u��[}�X��¥Ԛcjuew0��3�ja���E/����C��c����s�~���{�;�%���k�!�^��<���!Sno��)x�e�,B[���ja���۲Նɪk*n���T�X����1lenͻ%�`&��.�
�VͩpEXv�͘5��/7�}�l�%�;{�q���!e�ir��#��3�i#>�#��(Sޛ҇��W�+�X2��"j��B�,�%AH+LUp�����;��(�������"TmY,��KC+^V;uul��Ի�n���w����Շ�����r_���C��\诫Sn�}��Z��Ǎ$7�?��y��g��!�{����vg�w�󋲎`H�@��t���c.s��������:�ё���K��*i�Mۙ{+h)��]��Ԫt��T��%��Z��6'�>�6�����;WQ��:/�*�~��+Bg@�i�kԊ�{�ڤvt^,쭃������ٽO/0�04˱/9���%H���
ѷ���jҧ=���$ݩ"q)��0����=q�#�(q��f�(��0B� 2/9��Z�@TYp,z~+�E�/8ܐC�(s���NE��:��ͬ:�`�N@4�v�p]��
Ԅ�%8��m���'�G�<�j����یa��#���h��W�� �z�x��3�S㽾��w�1!A�j����$��:���K�=�D����¹���3��,񉃕N:N�}��O
�d0�;.��Ka�B�C�"[R�o��B-J��'��o@�r,��o��s�7�Ô-Q�jt��/���c3�1��s#�j�{������ ��:�`Jl�r�A6�N1s}^W�o�*��䉣/�p)��@ruڃ��<T�?t��:��w�SO{�y��l��,�ʥ�j�L�}.J��k��/�������ڔ��b=8�{�� P��z�����c�X5������ݾx@��g)��KwԿ��ӷ'�"���θ
m������G������[�|��&�5Շ�c�<o�1������d�3�׼���;��ŉR/�_+i�y�3Q��V��솒�~������`0��UmZ^S�T-#f��9e�3zG�� [�A�ڷ�G���V���*lʆ�z&L�냶�v��t��ݫ�:�6>���6�D�:��d�xF4�C6>:v�"�1Z��j���@X|-�� %�~�7��H��&f��x���Z�K���(�]F]:�򌢺��w^�Z�;��%ݪXN��٪mT��-ۣ�h��.��
�r��1��:��I�Y�c�e5���v���$kb�}y�q�Ɖ1�v�L��r��p�|�s,on������0'uo"m���@���< O1��b}�(��b��Rg�Z鸡����S
���6B��q�Mȓ�<!O8A �DqJ�kyYW5v�3���ؚ��NQV��2;�(����>�ټ9�.yX0�]��cH�s?%NT��Ek�Q��`VH�چ,2No�/X6���j��>�,z�t�z}��.n��n�^�=����PJ������[��t���IP�@b�RA�R�r�6�ڍ>��{���>�����83NO����ʅ�7@T
�4*9[z_��Ul�Rɵ"�0e�{J�[󒜳fG�<��VZ�|ɱL����C��|�g�I�x�0�plt�>����}�K�Rp�"G�Ksw��3m���~~=9\vj^7����8\�z���	��5���=�CY��롵�G�<4�=G�.7bl�I(5��4��zK�.a���LD�\��K�F��_/�,��tuE�%�)4��Yĩ�����ߢߓ�!1	�ۿ׹�x����*����k�E����`h�Vq���OF3��u�]�Qec��>Q�����Y��߷U���3��#������C��R��im����u�s�YV?>0��p�>�,�
UVWap��=lk�Ya�^�������˨0��@x��¸�bd���35V)�Kv�Yg�یT[[�����}����᫘�4�l���[���8QKM+\�0y��fЮ.Kk��E�u����߆q����=��%tY���R�2W_�sw(p�ڸS.k���M�-q1
q��!g�]��ƫ�))%����nC/�[X>�������f��Ɯ�+ه����v�/ɔ���1�ٜE�Wo@2g@�y!>�F�J��9�ܒ�(�`��ݦ���������d��ۉ
��U�q<�p#v�}�Ǿl���{C+�n^�使g��!��aE�t��-YlbKπ��J��lz"GڦF��z{�&|@�W"���C/2p��a���(��#Mk�ōX��,�z�.�TT��3��X���Ԉ�}+4V�3�56A=��5���Z����QÙ���ܷf�IM5��c�f�6���T�k��!���zG�zb��xU+�{�=�✻D5ŉ�K�6��Ά�3�>7��K��m�-�T'���.��H\Gj��Ϗ^oØ��7&jj0�����D���4?��4��X����'x�ݲKr����5�bRZ����gX'�m32hӤ��e=�a�y3#�`��N�v2Þ_@�������H�%���x�2�s9~���:U�AF�x^����G�1����(<���&�O5ٌ����=2Pm
Mp��8`�����ec䀻ǟ2���)v�d���:�ׇ4h�1��X {���kI�����ɯz�t��
����<�%�����qf}�=�G���b����v��U!��g�9����Rcvd��R����V�]W�a���t�ap��xW���^ޖ���Rۉ��K�ځ�21x���&�~mcc��W.�bì{'�3��aϰ�飋�8<�/d�1��5��Z�V�`��$jg	Y0ה6�s����*ɟ�y�,��31��b��$��m����ǟ�bE�j��q-��Why۪�̖�e R�-a���2jPmɾ�z(�O���xp v�I��7�Ῑ��[�;g��Mm��Nr�<��Z�Hus_�H��uW�t��Q�(i�u�;	�ܽ,�b}8Y�D�k�Xmk	X�8+�X�b�*���*��GgM�"��Ŀ�@"-�u��L���GrckuI���侏�{IF�+Ǵ�5�1Qc��!�Б�	(O��� ���1Ο{�)�X�;�9�J"����w�zx���-r�n��?@��w��3~O�e��2�IE"�����+���t��zq��8�����X���~�����K�&��ʮ�C��<Gu9��}v��?���8Y�K�G����+���F5�}E6�'�R�qݪ����dЃ�W%�*Z�������Sg������|���?�X���c]Ϩ(m�m��˴��%]XFG�Ȳ/�r����������S
�XN#�����K�[�����I^Ώ�>�ȼ	�X���3T�N�����J�7�u�چ�u�"�l~������К �ǥ.�1G�o�u��=H��n`g^V��Ӑ���"na��Q���Ylٷo�Tį���VNz�i�۪U-���v/�_��fs�b��ɽ�h����ó����Jq��~��ki�;�l��7n8���ߗG�}f�}&}.��?�֨�9���6��	xB�I5��GlQ��+9^.O��j����5m$w.x��v�c��o��NЄ��r2�ﰪYF_~���^�X����A�������$�S��N��Z���o��}y� }��8���b��m��'*�q�Q�\"���)�vc��� ��ӑ'�'�p+��D���I+'�K2,�x�͘�!��	��|�\tM%���D�g6[J�V�ĎGl�����+Y|�ӓ�s9D� ���g�"���E��~��1tm�$��g�dw�m�ƪNtzEԧE����+��_�b0&��ei9�!��-v�)�D]z���X3�r��E�w`6�c��5�4!_�T���.����w�Y�����7���%�I��v�B-�÷?;�R_���	���ON8�1 (�B3l�������;�Z��F��2"w^3��ud�.�"��i�k��ꫪ�~��wY��!�y��������ޜ��M�9���R~��?�I7-�n�y�w��H˓g��[1	�?7��3��3��Q)������
��3��� �/���1���c��%4<F^�}��9��C����_!HS\��������;n�-m��hi�z�Afkğ(��R<��C��ɚY�ߓE��!����� ��R�����\�f�N�M��g�\!�8�O�q����ܫ��S�nL	i!���Y��P����٠��z��Lon��������)��1���1�c�H���|��o��H�v�Ԍ�~�)�\9��<�$�!�,��96n%8�������e� �Rz�Q#��.��l�kt�E\N�������?���Cey�{O@q��Ε&�����<q�����-����a��q��=�����LU {�ko��v����{�=9�ۗ��?�YRd�N-K�T����B:)x���p��o���E��"�%	fϟ���-�t���G�Q���Ѐ*�������S����*n��F���=��c�\��~��f�+��Ζ�Yl���>J����*8�:&8�6��ot������Y������o��V(pRA��m%��W�`HN��J2��@�KU='y��i��9��;I/�~y��w��z���XF��k�u5���_�K�����W_=��{G;>� v�@����9]�cC7q��`��0���x��Q��&*ܪ������jJ��{�[����*���8/�Bf��=���-��`�\I,��Y�I|�A����M�c����V�3�Ԁ���2V���jR���Ԑ����J	��G���)y 0:�߃��:�}#�=پ������qb��]�a�t��qC�\L����uK����iX��8��z��/�[`���YeҺ����Ƭ��%��Z�M��H佧�t[���[�#��v���y���%�Ij�r��u�/M���8������������p���l��[q�~�v�{@O}\'����ճ1.��o��^q9gPE�W� 7QO֤0�Q<ǬN������L� �\!>��٤Dѥ�F����5�
�_�rv��/�uk�p���J��=�{ �annȝ�<�ȳ���?~�Pq�s�4��U�Y_��ߔ���ڠ�t�[_Y=�?������	���4��`�oF�>Q�Ŋ�I��Q��Ʒ=�o�{Ή˱�����+r���滩"���%�?:O�O���G M������7-ң�x.I�/7���\�J3M*=�dN��u1��s\ j),��Z.���N��SJ�s�z�ۭ�4#jc�U�Q9����a�|dh��+<��w`�2���S�;�6��՗~Η;O�s�}#��v�ɑu��Y��āB�o�j�&�"-������9�P��`L���r���#)N�p?���W<�{�ͲD�*9�醁��6P�V�IY��vڶ*��ǡA�3 zv�7&vT�H�S�%�.jvO�{�y��P:ac��9/�e�M���p����#��g����ob� bȂ�[�٬#��S�;O�k�BkQh��*��s[ �I��.ɓ	(���*)�A�H7'Z�_� �k����0�a��p�ף�4ˊ����@$�*���7����� `i_���ɕo��4�1��4X̓���rjH��>��9K��s�`'����f~�� ��$���G����tN���w�a'/"Ia8��S����V�!�iO��n���:�,wk*.��el�	�� �7JHhի�ʬ������e#Cb�)~�3e^`����O��ä���%qI�)��[%���R� <��~@\���u�&��`f+ň65e+�D��-͊9���e[�5���b�Uc@^��4Ǽ׈�jc�Mv��;H�����͵�J��х�^3�V����Ϩ� �K㮕{����mt�0/{/�0~Q����JvY����}u��J��� �Z�p���«�ƻ
\�jM��u�@����������H)�pK��Y��l��~X��{���٩��n������@qEBe��2_#�Q贄��/����"`;	1��nޜ��[� ��[Xi���v���ѧ �C`�����������2A���e�*����і��ٶ�Py\1�
'H�ֶ�6���� X����P��qc�->]�Ȫ��T�Ũ���r ��<.(|�M��|�s���w7��fO���=���#�	v���~�!O�qZ3!M� 2�hR�����c�E	�V���%���$�TL���h�̤u��	"�
$&c�;�$�~R��d��)v⡢{�;�Z�@����������:K2����EE��W�P�B��b������=0�km�����S�.^P��fr)}�R�&H�ʤ�����~D.��q%J�^�5���^��щE���K6ɞpqȘy�T,�-������/��T�'O�_���xs����-����\��b.�5iƙ��b\\*
�m�h������v�d}+��vZ�e�#d��䢻��
�){��L��:�-b�l��߿����Lb�D�!z�l�R~"���{�������<��{�/Y�ɶ�hR��P�{w��A�H�Cr�n)`�RW�{�eRUYS~9q���aK�O�S@��1��.�ր��Y
�hz��9�;�C���#�F�� ^3|3d��!U��pY(_�;|��sqN�\������
t�)���F��]�_��I�X��4|����Ů���Cy�.�~%h�O�Y����7:�����k5}�(�.$��� ��8�iQQyAo���`)�M~����r�(s���{Cˬ�|P%�~_(U��*k�.�9�[<�<?���7�a��;1��b/z���?
Z�Ī��{�  �k����k�ju'����ٻ!�"�5S:;	R��[�-b����������_	'��S1���.\��%�;>�`c�+�`fg-PX�����G9{0P�E����͖�Ǝ���+$�>�_����G�pe-л���g�	��{�(9���tE�UbF�
Y�?tP�jo��C���E*oG�^��1C<)�@��0�� �W2%�����dj ������E�"=2�@WA�B� �7���.��GA�wTO|�:���Y�F�5b�3��#7�A�� �Kl�66�C���\�4Qt,�����ц��#��.0x=�u�4H�/-W��^�R�5ۢ��~�z��������&qw�s�(����?�s,�we>�=ê>֤n��P�C_��Zv��u�Y��۟���v�oVt��V�};}�Պ�	����I�=�<=��.&�`,x-��m�}Ԉ_�.��}�L~Q�2�(j�tD�+\����.���52N~��?Pm���׃�d��X���Wo[EAޮ%J*r�Ow&��sV<����f���a��PWR@,"T��vtŢ��z���G?�dU�q`ͅ��U���ҵ�I'G>�JȼF�N�n����d�W&����n�xD�K�C�O��qw?)*�BI^�ɍ]
�?�g�-@�`9�v�ۍ������:Kwn���W�A<9f�1w����>g��x��H�8{;U�}X�@���E�/>���o����V�k���DU�Ug"�%K�+�}]ED���U�~W���B�j-g�Ɒ��*B�t���3�"F��8���D����կ�|? u>��R[�֐��?iq��`*Ef�V��74�-����w�C��m�\�Ĝ(@�|�W�!;��="��p�G(�*��6��]�	�����~����W,��U��P�i�Y���|���������A�6�au"�DI<��\�3t1?�����}P�,���� l�2S�F\+�`��; \��ۀ��T�EѼ����ΩL}���I�z�7(<������D���r$FP��v�&yn+$�'�D�C����f����ީ&7����b�!7)tX�^�⪘�[�(��R��9_�\6ʩ6�%\��ץ�|�i�ƈc�$ζ(TL��Y?�O�s��;���XMkD�s4m�B{B���Kޞ�v�*�Юj���S�k����f1��Wu6wbx����;6�M�G"�T��6������l~	�=�t���D��6VӴ���Tά�_N�% �ݾVRb���N+r�t�I��u�da�wvy��|x}0.w�����=z[�!���a!{��? ����BeB�	���!�B�ƫ�Z�V#��j� ?�|�� �P��$Ue=��ό©ފ���N�<6'��qϯ:��,Yʒ��b���` �<i��
����p�D}���/E�� ^�f@�?�}A-��c�����z�9l���R�f�`Vc;9�E�G�k]��p���R�J��`@��.�쬑Ju��ȁm�9.�9I=z*Q�f5�W�z�5M�I.u�ZE ���M�Q;�.�k_����kQ���U�l1�H8;�;��#�)����#�@{���f���� �9Xz���.����֘��>��3�����e�K곁�1�s�8o�sY���7�r�E+�$��_��ӯ��ѧ������z3� ����ٲ��P//��R�����<u���H����7���e�v��|B�
�޲e|t�A��y��4�K��3�$��7(��;��n{ '4�_*�x8Pùo.�V�p�w7i@D��"t���,�BW�5g���.�w|����J�׍7D���R.`g7<`��]7�rF�B�ׁ�J�-��EV�U;��h-#u\����p/þ%��ZpH���y q)��e���qk}y�GO� �u]L��߱_\ء��Yd�<n�i����
lO�2&�b�)���A4������f��W��� �w�X!��4��rY��@n�1!�AW޶E�cE\�S\��e���A�N���Sk?�J*:�]��4��%vn��z�ŷ5W� �\�z�
sݗvC����t�L|�@ L�k��L��.��o��s)j�l�%:�46��zp+d嵼�Ţ�K(o�H�L�V�z&���[�Tǉ9
xѨ*���]�ʷhji�g��"����.@u�NYR��^lK��x�xlG�vVz1.no�cI�hE��v��\dYeY;������$���y��g�(�j���tU49g���*fg����q��gQ��C�s5�����}|ڴ�]�B��l�����x��ܕ�T��CeOY;`�̊��`����Hz�շ���\��ό�Ծ�� �!�.�H����?\<O�lM3bw�d]�<����Evw��74F$pj�w`� �M;��!l#��;E�k�U��>۾��R.������J�~���X�Z�U~~Z'��BwxN�iÝJ��l����V�)�ۯ�'2��'�q���\�{:��ZQ5[����s�M�^2$�k3]W���ɋ9���𼒵Ν�9Z�''�	*��K.�#ͻk8��,��t8���D���F�m�z���ƽ89މf�u	)�}/,*7 Ҭ.�6�:g}��w��S�ή{�А�x,���f����*�B��/�w���ZZR�v>�3�:*#T�u��;xK1�"�k��M�H�wZ�i����0�⤃FoP��p#3�
��|�L���:�l��%[�Ky%�냘��e��O�i귇�O�Dht�P�/~�3l��B.��RU.��~�řk�z��f֔Tu� w����<{����>��1z�g:ŋ�x[R�<4C����b`(8s:�H�;�@������ypG��5��X�6���k�1�|��k������m35�1|�e��˯Ky�ݍ6�`w��{td6o�'�}�fB�^R��Q,~�k��6�H)��l��?����v�A��*��g�s�b78���f��Љ*�m�Vժ'�����SZ��^S��WD�ƛ+WT�`��A@ ���6��u��w�M~л��a_�jpB�Y�� �ݏe��Z�0E^��7�@#کU�ϣ��ҿ_��*����_$'һ�r��}�~��M^P�C
^���P���"���J��\�^�૓e�+��B�f!�u�ޗ�eUt�M�7N�&�@�.�s�v�уD�{�[��ocB��#Î������c�2�q�ȃJ+d|]�����9�+wb����c��� ���M������Գ���sg�Qr,~}Sе/�g�+P�w�f�8���-�V��W\���~��J������n1�;2��\Y���T�+�t=�u5{iuX�����$s�%'��e2�q����۷*%��������}[2��M�Y�ڛ-�֓���0�w'�hR���,<��1ԋ ]2G7�<������F�������}֩w'	�����z���;i�qR.+���e~q�в͸c#�f@��Z�eq��f۱�+�������B
|ܠ�{�c�U��.\j�c���Ä��\��k6nQt�k#�ً?Fn�~��o���̘��^q�}��� �'��p�^�W+���4 ���h��͝!و
XNV(Z��蓟��~{'�'��ҷ,�v�"D�+Oغ��]��-t�D_R~�q�����Ph��N^r�_��-e�J�Uڢ��r�V�f����'�z#���7�@g_5��� XhKyHQϣB�9�Q~����i^�c�b=�J<>�p3�y��>����~ex�Eb|�+�_>���p����%@��?����~Qww9��\���3�� ��Vire틑���$ε�� ��3<��Ι�k��00�}�Y�]����[��4-\�
[��j���X��
1Vo�	�_�*�9F@���4�I��p���i�x���*5��g��Y�k��蝁o���5B�j�{�`�F����j���MjGE'WH�6+:��CO�F���`�&׊v�GU��@�������@��tiJ}�~o��IoIB^��Mp��f+�C>�3��ͨ!���J�h�m���K�cǑz����3��4s�����lE�Hu�f�md <�\A'�L��D����{w^M���g��-�P�֗	�ׁͣ��Ђ��ǂ���.5!~*Ë�'պ����q}�
 �7u�`E�M^�#:�n*��G��2�m��~R`5?ЫX�(�5��X�<����c�E�.���t1�&��,�d�`���k3��6�*����P��W=?�ƍ� KrZ�ؿ�����ؒ��I�r�q��»D���J�tM�b�<�j�mp0�~>�vXΫK��8aH�m�z$UN��~�{&um�2��Cr���1O��6pj����X"��o�ޯ,~R�;e� �l� ұ+���t�⢸�Y�EE��0es�qYVHw���L�n�KT*u���pԠ�:�&@�7&u!t���$��\[��Awm��_ܺ'�Py@ɸ����� �1��f���e]��_�(kR���n���FM����y`�~͛��}����|�F���޵��2��k�,�@>I�"��B�ǂk�#F�*)�bT�A{	��M�%�t���4�(��mG�-/��Jٗ}����D�wa���W�`�Uxb* �������*8w2ݟM�{����l^����$f�933����E�z��O�I��
j� ���5[6����+'���$�x�r�����qtzkmc�?�DuCf�&F^�sO�rk�s'O����oG�i_$��|��W��v=��遅�S3�FZ�9�d1!����0�U^(�"�UA�H>eS�H���<�tQL�|$KeZ#�T��e}M��J������i�I�x�C�cQ������P��!O��J2;�VSF�ٱ��ݜ��"q�[����� ��7~���4�نϷ}�O]���)
a�q�f�{6�Q<���y�����g��S�FnI����$4�	B�[nA���Ěl?�&�2S/J$�8�]�v��v��V���p �\T1���ў�4*:�vu2����0 F� ��Tp,��[S��`6o����buG�ؔ���$(Q�+l�*���M��Tu̶�G���'���k��*�0i�`%�F��#�D�x�0�gia�噐�֗+[�1��ئ���+�4�r�%ǥ*��	���_ȫ7&�5P��J��A1*~���I3e5�D�g�����lUߊ��dWζ����$������+��7��/m����r�e�����sy�m��]/�70�69e��t�O�9c��B�R�����jچ��mZ�P�/�o���Km+O�4Z���|*&c5�w�Z(��Uږ���<~�r��fN�p���`0����U�{��v�i���c������>���_!OZ{�(
I�Z]cQ���5���-v�:�����g�W���
�a�U�{�Nw�{^��e��aMsJ�s����ӊu���c�~\s�yJ�g���&����K�2�&�zEH5):RǷH��K^�>�P�����~B}\���D� �� �����7�N��}_�oo}��$��V�+JJ���z7i;��I��j��-"x~�|-���HgbnvT-ǲ��(dK{�F��o?{)@QL��\�]�]9H��'mz�+sk8�j�%qE��Ee`���K�RڔF�5g��(mu퇹F��i�-���v�o�yq��-AF�r�3s�E��9ɪek��g�SY�,s[#�*�����l4ٺ_�$N�4�c)K��f�CF�/��"��
�6�4�W��+��(<:����u�&��I]�Ď��0k�}$=���/����C-�4�7��k�P���`8��8"E���)�@�qY/c��>�{A,?���f���4"dǼ�o�������l��G�������?`F��^�Zyum�O4ױf�'�,����~�wCUG�n�Z�K��K�~��+�YhQx���D�8#|Z����cLK�����o�K����j�]6Z�F�S�G��V�c֝Ȥ�WQ�'24Q��rKԷ$Mθ���╗�C�jS؋âق����v���cv�~+�0�}v�gE;��t9g=��is����<�)����2`�fy\����|nU<��_H��	:�\H Z(Y�$a}�!�c�0�Q-E����W�$�:��`AE�+q
�|���:*�{sb��Zxf�Rr��/\d�
���7E)��1�@���.T�Wa#3qp��&8�������E�&�%P�b}i�5����rη�N�	����h��3��>j�^�\��wB܅�S=���W$n=��1;�r�w�v���M=��e�:���Ҳ}u�Tq�_�F�_Sj��dٽ�Y �?J�'��=�1D�}��{f�z��"�������k�f��s�ר魵1�j�j�� ��P59��m�D:�3�@���q8N�w�� WA�?@��	�'0=~���މ�|ڭ)���
��v=�@Y̖����Nn�ƱꐑZ?#P\��	�jj@�'*�ݑ6�غnW���Z-D��	$�������]��݋�Cr#�T�{؃�߮�yX�y/�a~���A����)ٸ��3#����-�a'԰,�)���1�K�n��r��4Ɋ�N��@�'n���b�E�aU�������5�"&R3�H�z�yᩎ�V�soO��<��8��>W���$�q�pn�룔�����"&0J%�˱Y�����>�Qq�r�.3������nD��`��$+M�7#���"3�B�xV���HbǞU������|��_�yա>�c�@h�����_Y}�ݻ�A�]_���H���Uh*`wN��:z���롃<��}\�f|���ve������C�7&����_����EU��xCС�J�Lm���+���`�/�
��2����k6[��;�v��.���{�#��֪�h��K�Jճ�[l��u���[�2/|�9�^��/��9]�W�+@變 &&���o�ĖU�h�Cј�5����l���1j��W��A*o�'�w��T���")&]O ��bm����[_H"����b����lq�ܕ�J��@�Ow3p/l`�!'��aW�����XX����x'h������?�Y$�X��ɫ����v��%�y�z�Ԕ���D�a�e=��4wW���O�e<�]/�h�|���2ooƿiZ:>�m���pN�+c��-/V�	6
^���͵l#jA ���$�z�8")�+�i�r1Z-����
�cB�&a�6��fu�߼<ԴUO����]�KO�4';�&�,��\r��'J!*_����Ư>�ne���MV!�D�*�XH2�vo�V����a������M-G��:��.>�lH��z��o�[�X��=���c��ܧ��M��]P9_p5?m9&<�(�jv�J�҈P<���㳝oqk[/�nLte���|�k���i��f�jI��6�X�Ja�gw������͐ �ӏ+A��U��<V�Pg�XLupO~'Dc9\�k{X�2m����(Oyq�,��6�7Dbk��험 �b��~�$v�Q�)�S��+��PA$�	��Y ����&�Α�oOl��7d�_̩�f�;�I���G;n�}G�ˏk#���W��A¸���:�A�c,�`�����;! ��F��G�}}��h���A��î�Q�\�B�i���Ogf����vn���렟�t�����M��e}���F�k�}�8����ҝ�]�iAZ�{t#���������������b��8��y}o�v��wg�tj%�{�_���O��3._i�L�[���Q&��[Gz�be�MX�/3y�P�s��e����;%��7�@��fIs�,���>_h)�:ʃcĐS����>�Y��l��c��nlJ��D��� ��UYIw�̂�����L�C$�v- �ȳ��"�2e#3��4%�IwQq�� 3yX��Z��D�$g����p��.������n1o�z]ht����n����/�7&cN����Y��%q��2��9���r׶B�	e�9@��E8�(O�+��0���K����m��#�m�����l������S�X�z���q/�
�:�4�j���H|����I�Ϲǖ��̭7��E�hTr,�PZ�I�@�͆�2�q�G`��߮�[f�������:�f)(?�������P��t4]d��p0Xv�ѣ�Y�Ө]�9of,i�٣1��ʾF�/0t�^J��w+�m�1�ʬ���,����Ԫ�Ȳ��=ʕu}.�ؼ��>ڐ�t`�"%����X��X�Y+����$2,�2�`O�thN���-Y�,o-���_�	8����l3]���*��CQ�%L��H::����ͥ}Y�Շ����	|'�����kq��C�pW��s�����eJ���o�@0"	�g�cɫ����._L҃3���}��,,,�����v���R�g�\���=�zL��5ɲIΥ���gW˒�VR<S�g�Օ{��o�s.�b��<M)F���e$̭�c�hЫC	��u1�<N�0�G��!�M����N>�i8i0[ϨG��j),^9)L֙����^`���Ե
'ݏ�F�C9��mKf�i����B�/�[�;f��_�hC3c2�.��tC��ǝ�4�3������0�\[�ˍ�/O}��e�����;�.��Z^�v�u����4��G�AY��n�7-l��=c�n�T�Dc6�w�Xߋ�~���@���m��@��$r�|��>*�Q�2u��ҳ���(�9�#�?��-g�I�z�C�2b�C�~91��-��k��n]{�x������{9lT�Ջ�ϐ���r���Hð6QS��g'�����ٺ�>��U/�$�;�J�!�ɘ��}󄞫�{9��w���p�<7��-���a��!��R���Jd��I�a����<e� �AK��!�R�y��k��e��#�Ͼ��sT��u�p�	�=�iz�:�#�s̸k��&)R9�^}c�J������;XyX��;��Wa�#͸U�V�u+z��G����| �3�j$_B��Ջ�@�:,v��X��Q/��@��Eފ��L��)Ί^��RF3�U�����Og����lg�'R��j�A�mj*×y��S�d���@�:�^=�'�ٷ1V�⒕a���E�����ҍ��;.[���������7'խ]��;N�ۚ�<*F�p~�}YHd���u�@:--g��;���������扆�i��Z)��#;��{?����>�%��4����<L ?�di�ޭ�	؁ڌԧ	�����U�Q�^}~6�'���{ڜ��	|����y�d��A�f�6+�\O&n���ܾ�:��p�}[=ֽy��b-�&9�Q�0ǅ�>+^g�6��\�yy	S�XB�����nN~S/*���D���O����ox���q� ��^�*��Oٽ=Is�M�>��4����.]x��]��YRY��I*=M��G������z�\�e&K?u���
�/^[W�n����b�k}군�*���R�c���NI��&o����C�וY��к8���a�� ^ן�C�$��c��`ħ��$�ٚ����.1L�v ��c��^���:�����lh��m����̛�^��Jǅ8) *��ᒅ����^�|�]�{!�v;·��Ƙ�?��g�����%'h���v�A��� ��	}9L�hu�@#�ƿ٤���>��f�\����w6�n�F_!���	�Sܸ'��<TǮ���Dߣ�׉�rp�қ����^���ޡڴӌ�#>����u�I�D��~������S֎����N6����jl !يB��e�-��{��럃v�I�C$*�����
�m}T��Q�ә~����MEsɔ�;zn������٤Aw�âe�ңu�1r�C'������}�XƇ~�yvGx'��w~�%�Ҵ��8�V�;�|��CGq�c�x��2���/��`�׋��{i�p9��Źn��W�t����N,�k�#�}�R�=i�o�R��p�7��̖��k����m�-��5q��ҭO ��;���{s�ýF|(���洭N-�����l�_���!��
���e�W����N�`�v��X6���G24�6]3�R%UP�
�3�O|k�*4wWP�H��C��4`7��$����OX71	���z��.I����uw媵��W�	�����"L5sn���H:>HNZ;��.Y[��:s��NJw����v��f"����߯ŵ��������׫�>���� 4�~[��;Deo���>�Ʒ$tAHȢ�E�[���W]r�� ݀.���Js9mfˬ#��
)f��HoD�57Hgz�� ���o��D��g��z�*�H ������6|	�x��
=�U�K���olQNq��Yϥe���b����̄���7����Q�'-IE�f��_���Q�Ѽ����ϛ���Q��ዞ�wS�~�{���Պ�u=�=R�<�چ��og�B�@_g�"Ӧ:�u.*dg?ŝ<d[s�d V�E��J8nx�4�,aoڿ�z;�Ǥ!<J�'��A۽�0��n���
��$5�Ook��1��&Һ��<O(Z���Yt�i}�5H���t����-OV^�w\|ymF�a�e��4&�F�~�v���| iV�8*�Le�*�v�5<X�V���-`b�͓u�����Kp��E�l�v/��CQ�ٮ��L���L�}|smB90IS:�x��$�ɑo�y$lwU���^��&j�q�$|ȃ�f�N{�L�uJ��ޱ(�3ˀe�$�ck�&ˑ�ٖδqh^�"d$|��4,Lm�#��b�wJ������p+~�.
>~���d�?�Ŵպ���A�S	��#4�r\�3�ZNA�|=q;��&��h��{�]{C��i\|���ݐ}%�αx
���n���lC�0֊��e�س�����T���H�,��
1�Y����e�c�گ#��u,_W�67����'��@����+����-��%^��eF?�*C@��ɪF�3��*T�.��φ٦v3�[�?p�[њ�Æ����^��2gDG�.��c$X,�ƅ��:5�k仇޹l��{�%�3���i�>8�$�����Dv��B���VJPh�'�S(���*xJPϖ�k��I����h��|�OV�"��L2ۊv�*�M{�4��7A`W���5��k@H`>}486�D���M�	�GIJm��~"k�u6����a���ay��?)�����
2�pg~��>�?p���,v�-$��2>y�MBA����R`z�P�q�h^�/.����<)������|^qxr�y����drR��i���f(�~/x�V?%��=�W*��:VL��@����N�d8A���L#��χr)�pyvM`��o.�rf�0�������Ҕ f�����H���$��+�"T=��.,�Zd���k)�%J�Ǖ
�B�(�ӪPO-�\n̏����CRs8�_ɟ��2�?n7�&�Y�Vm-��ϣ2V��(h��P�
s�<�����}{��%o��(�%��'V��Se���d��@�����8���*U(	�c%�^z�ya��2�^Y> �j�u�jѧ�$����ruF�5�������<Z"U��,[~���o0�1ʪl<�?�e>��8�m�NO+��R<~�d^�I���~�����^=��Sȯ�� �s�]oSU��Տ�q^�m��(!� 8sNN�e���ܜB���ܳ���S
��c-a'wF	���+���<0��ZE*O�z,���8�-�0u���f3C�*;x_��'�8��WQ�z�����U�i7oqv�[��,�է�{L�ܡ���DrH�#?&���Ա����D�u�!�,3�r̳�"!�SkF$�g��"E�DV0je���]T�_ĐX�
~�ڢxd��6U���HIg�O����G*5O*'	-���gl�Eth ^�K�����
�g���8 �˖�5|�"]��9�p��X�[�H���L�n�-[�:�+�ӷ�^�_rC��F5� ���^��G7�W,8�63��MBY5�7S�<�Q�A*��TO(Գ%by����粭v�'�a+���>ߏ}�}����ɳ
N#A�O�Y��'g��#!m�%
ܑ���`�TB� f���^�4�W�_�O���2���ZIe�2�[?�����'�(�DX�!��G�k�8;wda������]u[�_Zb����̤D�:��X(�Q�kcQhS�~����3���O0��pwDXٲ�[ ���{b�G	�6�3 9b�e�#�������ݯeM�ۼM�K �O���x�D@��J�B���J@��dm��C�X����Yƌ�O��~�ڽ��+�u���0 '�1�U���{s�SA�����n��;���>?�L0�%������Is�$t�˾Ok�� �ڮ�*$Z'�?���ݮ���.����l��P�T�͓\�Y������W,�Pc.w8���*Ux~��ڱ��dd�Rd8�_�=��P�-#����WP��H��G�ث�y���L6�!��de��|8���9���G�����:^w)�\�?,L���kV� ���PQ>�c���>d�	eu���}[ZB=͛�]}��֭
��M�	"�<mXB �����O�f u{���
��6�[衮U�7�n��/d����	��*�8����Y�)nw��)ۀ�ٝϵ�>+��~��߰v�a�|ʞ���������"����|�ha�S���?\���}��~�<zٗd��{s>�U^�E��3�s ����,{�#_\8��dk]go܄��a����3#���e�a�<�����}�d��Ϭt�	�P����0�W��.�qe*��.�J��Z�ˆ�枣�i���	�����M}3�@����B�48���{S�vl�.�
Kov��-�':��蜁����"�8���zv+h�6-4@�߰����1:_ŀ�
�nqü�f �}V:�q���]r��:�쁒P Ժ��Y3?�]@��ӵA>5�mm����]+��W��!����|��W�n�ܔ7����#PK:6Q��/B^��kz����S	,3�f����T��l���i��="[��-��4�:L&�rb;��$ᜢE\V�n�'��/�0�!�r	��ob�zÓ����g}���/��Q�Q�RcovWG����a����@�Up[=Zê��
��u�A�i��6�X�C��x{?i�$�D�s���,u���6�huZ�
9�����5Ϗ	ӑ�E|��چ1~g�st�ˆ���!����a/���������L�/���.	R�E��*ݒ^Rd=Ѽ~�ghma����,91t;��\�>N~�n�YA���&il�,n�v���R��ϿnT�w�Y<�/�������?6��5��S�d���"��1���4�I�8�S�E-�p�SyT���H�Z��W���(��ۙ,��7כ�֙��.��:N��kC��C�p�'2M�T"�}ԁ�"e5�]�;&�MiB��.o��I9饽�,���&m;�g]G�t{C8����[w}$^�k���侰z�(�������X�`�C��`��j�ʏ ��O��VJ6�@s���M6i�3�5��"z�=���9�e�Z�P���r���P��]�+׊>z���c=P쏛��c�})u�������C&5R�ڼV�PQ�N�����3ԉ����6����G2(�l&�s���������[�l���w��2�[��H+؄�A�U��]���;+vU��)bGy�����ޜ���:���� ��4�ä>�u?ڞ����-���:����ޫ�k{퉺W	W����{�.�ϓQ�U�>�D�à�Qq�j����g��nx_��ci�ݙ�I?���`���pF� �������犓U�19U�Zӽ�uJz����[H�u���3���N�88���!&�ůr�p���d Xz��!m�j�p�]���r�|~sSwvX3�x���
n�tJ�跖��x�t�82�=zE|�%(�@�O��d����WoR}�K�݀�������A-ϔ���$R��9T�z�B�rG�0_j'�pa"�倉�7ȹD�@XO��.K�5�����~�pTAj�'�_�s�~��A�}Y� mh_�/Ɍ6 �=h�b%	Ɇk���E��q'�il�}T"Y�p{�k��t����;m�>M�z�'�-�Z&�f?u';<�M+���<1�q�����
��4���q�m���i��WK����B
�l�ԑe1�w(@jZ���9���ξ9�\2���\�FN?��
܊������?��`�A	�i��ځ����,���Uu�Oy��ql����)Y4�wK����=��^E:�1�>P����x8?ZX5�^���4��W8�U��4�ډ���H�$?�&���S�����9`�ON��=�p�݊ ��ޭ��`�����콩��������Z<��&2�g7_
^7�ߕ�>��"�^t`�x/e?��t�q���� �x".*y�C{�Z퍪KpB�Ex�C0��F��3|pz��R�=T$��uvZ�U�������} w�ҟ�����0�u��a��~��<��]�A�9��{���Yk���V����A��*#���%lʤ���B���6�]�!�:-�X �̇t�&P������~��#T�r��$x;�D��	��5������n'￿�&��V���$D��	CMp����b�`����^Ӣva2w�]P%�S�wQ�|A�&A^h�V-�M^ ��B������?���qLҕoV�������)�c�*��������D�g��n��l�0I�0�$�����E���tA��7o�n's��j7Og��A�Uo�&I�Z&�o�Ӕ��%� �e>q^����wr�m��c��/k#ݨ�5Je��٣�'|-A���
��60��` ��|�b�H''�9�|T���n��σ�/xCV�%�({�����\���-Ҫ�T5DՇ��ն�'�f�������=��a�L��?��RU-P�*r��n�+4�zQ:�M���x�>�>�����D�aI�ߗ���N�O��㾆��?�7�:-�9�::�L\��p�7�ֺ����X�u?b����p��O/;y$gkW=Y�K���#���"G[x0~,
�<����S}y ʬ��Ϥ��+_w��8f��2�L��AKj�9��<�B|v`�P�n���.y%pCT5�O<NS}��@�|!ǘf�z��G��G-:��la�?Z���r:�9z���!��4F�벬=u7˴���gemOX�8ǧ��בM�=�z�Z���=Aϣ%{�J֮�Q?43��Z�eF�`���mE��D�R9���[�p�6�q�b9�7��ma[��o�ǚ�׈q�ű(�]1���C�8.��/�u�d�
0��S�����͗����x��x�Z�����<um��w�����Ȭ�-�C3=Mi��cW�Wp�8�CF�Ҝ��[��φ:�����_\dTV��?-;}��{@�������0%㝦hɲ�[2 ��#��6��=�C���X4���^N1�pc=]���>
�C�����{�6�k�8�vI�5O,�1S�B�~��0�#�5�F�Fg]M���R�{�h�8K��H���ГӶW�c�7ڷ�����߮��2��3�D���l���3ƌ�bn��ܟv���aܽ�����a����`�z��dE�x����U
ɽ����1��u^��mo���"��܏��-���9C�ij��(��-�"�K=�ҽ���y�R5N_(vvi�*��j¯uA�k��h[{_�g���J�w�g���>B>'���N:��`�*�zR�D��4m�[w��¦߬����<\�eެ��rst����?"�������1��o�_�K�DT�4��a}h�`H�O��6���Nf��u �%�ߕܵ(����f�	���J��L�q�nzq?Bu����uڻT�6~���{D8�#۽�&��%^&��p�VX��<8��0IcN�Cc��B7��Kk������2�lr� C'ym.k�(S�B�%����E�Ԗ��l��h��R٤��ș��p�u�]�n��<��<j�ҊU�N{�^-�5T���Ź*�P���w�]G�������z�7�5;�~��sia{Q'_U��~q\y1����K�-��2���D�o�p�?������n]-����W1��@RX�wS��1ɀ�T��x�f\D8��.s�&$߬ )��ȓ��.k�aK֩�hё{n����h��bN���oMr܇���,�,�XNCT�p_�k}����Uɬʡ�k�̊��L"�ח�>�i�4f�����l����<[���e��w)�+|��s6#/Uq���V:������%���83~f%,[Q��R<��ې�&	9��T�Ƣ�%] L9�秌VMU�.P���>��,�Ζ��d�WC5G�7�Zţ
mli�waM"E�m��8˹8���'yf7g��6ZP Gxt�z?�ְ��y�2O��kko�io��4 f�}S�V81A��^�����:��4���yP�|�HA4^�����'n����7H[�E���O�Qju�Qg�r��齱;^��z��˞ɷXj"z|zq|w�I�V��z��CB~�節�;+I��96�b��J#����q�F&��eY�q��h���}�'4g�2����礣<7H㫳~UI�+~�*��m�쎗iq{h��)��Gn
��]"�!����Ԧy�o<��ӕ�ۣO4\&3_�
�VE����*�����>2ߢ����.����0Re�@�y��F��ۑ❭��ܣ�s��\��76Hk����¨j�P�6,s�h1�3{(\�n6�v^�k��}��A杓|"�"��]�AI�	���l͗^ͼP���M��C���p"-]�D����F�)%��8B6��!�%��]Ϝ��8����E�;���j�m�2MI�/���{��,��B�Ƙ�&��)�(�^ΚK^^Y��_�#,us{|�]4�|��)U<� �Kj~%��IF��4�t [��2��VE���(��Yv��~�|��u�I-ipr��ԧ�w6�Y#�[qbfjyr�����в�+*�#*QǢߺn�\t!ץ��u��/��W`!�l�n?�ʬ�GÁ�����k����ZuA�ʳ��@Ȟ�k��K�\F�ڐ�|d{�Ⱦ��3|P�2Z��YqP=#SZ��Gg�{�����_��҄JB+����=�n8靧V�5�v��Lu9󖿑���� ���!���gWw�l��abPS*����k����_2�6���Tg��Ɛ��q��̱�J�ş�Uݓ�{�h��Mx7��4΋{i�fFz�ǚ�1lh�S3��Y��e�A���=U�E-��Y�����
Sj��;��0�cCǷ��kD��<UB���{{W�\���Z��;�I��r}P�grʊV���8�k��6N���wי���\��׋��wf�����\~dK�]�5V����|�_�G:NW��B{��?��6��d��ڊ�.�槚�Q�������v�䈪�s���B�O ��gz�'���*=}կ�!���m��8?;D�7<��>�']!�����U?5.OQR`��>�_L�>3�R����
.�o񘑘�=B�WE/�x�:���v���7^�<�M�����@�u�-B:��K����A^��ff���, mx~��ۿ�x��������C������
�o�# �e����K
؂�%c_�Y1�+3w�	��B�&go�J�gLo�6)�`gC������a'b���x�E{�?]5��3�Y�QRp�����J������a0r�����xPpyg��dsy�.G�^�?�F˅��S�?� ��|ZN����z���U4�p���F���'����o[)�����p� �l��j�;�+���P	�q��+p����߇I(Ar��%0��YH�mQÌ��T��ΨㆸΨ�o����;���Q�� ����r2 `�r�c�����q����P�K�s�I����V�ݘ�|��;o�kh��K�9��x��񰯦���s�_现���n�C�DO���B���ԟ�^S!O�n�N̰ho�O��6�I����h�\f�;,Gw����B���>�.���2_6��UHӬ��.ֹ���Omi�����̾`z�ed�8)��]�l;s��Q���3 �.(�����]z�:��@ݝ�������
�q"���[Z���fo,����/��.E.z�=ˁw�7��S�7���-����j�����DQ��1���iIkW�L�4�P�sp�5˩��"/��Uv����o��\�99��,�������i��FK�Wx#�9�AGVV.(W/�+7ڻ��l%T�	�(��NBL�C��xЋ�j��yL\�p[Uj��.F!��?��jʢi�^�#��*�$� v����'ۛYN�VF���~����4Btx/v��J��������r'�d3�طb���e�dK%��Cw��Y��2�<LNY��b3�4��֒U���S�*��g�-,�Fi@#��l��%����JԷ�_��Uգ���)�d�wr*�5�5I.*�p-ӓ��Ǭ��Σ	��R�]�I]?���MW�ؗ�,�ɬc
C7c�����&�	X���l�u��k��6��|<{�^��d"RItf�-�X;i����'��'6���G{xꊲ��p����"�[�����N,�� �]���O��
��q�z~�ÜN'o�/5ԩ���Ǘ��P�%�{��/���X�b�T><�/�~��=s �5�c!�B�O�L��f�aS������`+x���vf�<��[98������GW���6Nm$�.�-<�Pe�V485�W�o��(�<?=w�|�h߱��œ,�c?����|2;fｋ!��)F�A�N����	u�O�j��A����'Qi��i1�ߦ�%�v���A��"?�	`�JOx��ҏbQ���g���2�"�u�f'�m*���2�)k���6f�H�/܉@����ԛ�ܻ�ʌ
K޺���S?~b��n��f���;4�H��o%/��*���k�QT��/u���v3���p����r]�a9�1�cB�]���zu��	ޫIF�©#2�(���R���r�)Ԗͷ��:��}��cy���Y�)q(+��+��Y���[dȴ%�,Z�~���u���[���R4
D�xy�+�|���?��f��Ĥ���/Q4�i�=z|�7��*/���.���ug��Z6��CЃUM�xݟ��oA_R�u������M�� 2�mW�z�,
��k��5�1��?�����J�n���ڂ�W{�k�ž��}/�n�']Ԣ9���۵�l�p�*����#C!_�qoiw���TpB0�)�ٹѫ$�s>�#7e�}�ڷ�f���$��������W8l70��e)�ß~|��1��N�����$G�ܽ���+Tk!3�!~����'{��"n�,!�W���h�<���ސ,��M�@o���0���:�j��&7! �$R�ke�ͽ�@���!�H��r�ݿ���h�-_��-�j�)pվ�*F֊p�F�`u�v�$?��m[��~ٜE�RB;N�D#�F�@�;���i[�Jӽ��5��oG��ĞykV�L�����|A|�}�7��fb<�o��vG
Gڨ}E�0uY��C�88��jCHO3���ſg�a���}[�����n����۲�SɎ16g[���$˅�;c�y��0��Y��X�GDkA�\Y4�Z�Y����B�W;���*��Q'*�F�w��=�ϔͯ�5�O�p�4lF%�b�e~���T�H����8c�䎲R��܉����^3�����^vk>������;;�x����+iOa�f.|t�H����S��ytˇn��E	�����M����Ux>H|(�O�P&w�0xW7��Aȯ%���akm%��:��ʻ�0��7���5ot��(ܥ�����R��Z�/5�̄�^��A{R�F���d���t�$h�i������ݜ���p��k�56�n����~��Z:ߋr�%�S�m��ClO�w����N()h�#7p�V�4Dk���/�Q��C� )��_��ـ�����b�\�E���l 鏙dDA�E��J�<�*�5���C��;
�"��2��¢Oq�K�{��3{�X�y�.P���������~L��*�E%��Pi�o?����h8��u)~�b6z����,M��]�Ÿy��흙�H�7 vEV��6��uE9��y�.��=�9"A+�}R�<P���ď�sSqy�����X*=K�������ɺmP�:���o��s���s��0_RIf������^�d'�}I�8M��Ne9L�T�k-"�;Aɲ:��d��W�|8j`P�S%Σ�	�qK����/��bv�A��
�J➣�d򑿍�)��*fU E�&��Jn,:��-Ol����=
��mgx5���ě�4iȲ�JC��?6�wΚ�c��k+�D_�g�t�����n�&�-o
ͻ+�����w�2d�0�aà�c�Oܮ���F�U�o_���?C�����:�Ӝ[�;)P!�W`���u���� �I�`u4_�ڰ�t�l�ȯ��6��<�R� B3�h����!����U� �x�?1��qȭ;:�Tн�IV��Ԝ����['�����tU��?���becs�0_���{��Wf8��'o�LB�7W���?T�)�is��'��v����xB��شxu�-��]��S��Β�W�`�b{w��	��Wx���^p�4�4��$��2b�ܱt�l7S%� ��+B���N٥���ȡc/�A)�Ydc�,��"����q�ç"���&��X��M��̚��a�m�;IWK�ixO��&-��8�ϊ�DD���P���m:`�3��ғ�t��@[7\4�a���B��O"=N="�D��Em��r���F�m�ڱ���+�R�t���4�ԓ
�@�N�ܮ'�=y�������?D���hv����w���*^��l��BQ��ְ����s��F��%�x�eX�R�lڇB5L���g��n�jF2���:�2LFKyJ����7m1n��
w�k�D�8�DȾ�5|�z屹����?#���]8��(�#U�9/���K�R��bY(n�����Ter�9Q&Xn����pk�lk����bHd�C�}8��c�mrvk�l�0dL�&���ʗ�:��i��?�{m2�G�F/F���z?��gƱ��-l��ݥ����~{?��7U��D��W��꼮6���)�$��&�)�����Vq�.����3.�K�k�̩%$R����J���x ?Ie��\������~l��$%�&�R'��l�9[�L�6&�� ҃�Q��{bl��X��X&�i���#k2��e";2	xzl�8����֩j4U�@��(Z�����4tnA�M���[u,�ŋ}���9�^G$Jː�kϪ����{�� �:�6�����qvś���7!�c��{���[!�G��}�	�O�������n�_TA?� ��w���?�?%%�ރN��M��2��	t�i���	����f�vX�����W0x#y�O�u:T3�ۙP�
U��\_����l$���#���x���i��ka��iQ�p�&������O�'v��I�Wn��"5�|ӿ���tȫ���M����o��U@?��jݷJו��[]�H�P�U$`.�m�lB�#��f�be2�}���z^ ;������&��\*�][�ъ�ֽ�zi��Oֺ+27�N��C���A�W����c��Zbd"�ȭ����n~"S��[R̽o�!8�b�\�� �	��j��P�~E9v��54)�ciy�a�*+���+N�k�˓sߝ+>��K�����l��t^K�h\{7���/-Yl�G��0Q�����D&zj�.I&�|Ȍ��&_s��ݞ��4 ޴��
_h��,�����}V(r�ڔ[�>`��蔆���A>zk���0n�_(�ْ�m�Q�q{���Eof��g�t�Ը����oe̓�>��UAC^�27�҂Ŧ�oȰ�h�|�{f[�H�=yx�j[[TkY�=�-�X˗�IR��ѫ�Y�[T]#<�"��>��H������W�� ���\{j���kΈ-��c1 �SX����+\��FE̜�ǻ�~=���t
L/�w�gaW�v�Ce4��A�S����W�������3=e���ˇ����y���Q�8�W��/��P���'��c Q�lQ�o�D���ψ`x��_�!�@jWC�W�y���Aщ�g�<#Ҹ�t"VW7Z�	�΁��蠖�����2Z���H��H�Cw��Mo��f�n^R]A����v�����.��F@��fU�~ٚ�,��V���`��������rV�ԑ  �{�'��i�\���W�!-<���0�O��v*�����g1�kIɆ ��� 4UȖ��u�~�5fL��y��i�2��p��{J��פ���������hH��0�2c��[el]�b�x.Ư_N~>-pP��ƕ����[N�Y���"��-�*�VC�O:b�^'E6�7���9�J��*�z������`;��5v�Mgj�����lk�2<-%����i�Or�������Wg�M�r�����"�B����H���i �Nh�����!V���	㴆8̐���⌤�־�G59�JK�3���;�4�2jc���YÐr��2���R��n�����R%���E�Ǒ9�X���aYd��b�?�`A��^��0[�ǈ�a�6.I���eGѫ�M���5��W"�&�Y7�ήl��K��A�]���E2��2d�Y����3ZI#oPE�F`���#x�%�Խ!���E��4�V/�Tfބ�G�a��٥���m�p�S�h)�Im#Cz�2�C�*�"�M}A!����;�Q��o�8��޶0�(��+��>�l�Oئ4h��ʻ�� [)i\[:'���m�l�u�xQ�����#bqBS&qq�پ�W�u}��
/_\A.��_մ!M�bn|��f�����u���~���ĲT�I�������7��Q�}�v)3*K�&�5�ކ|��;���X)��k�-����3���m0�d,�uW٫0�)���!��hF���c͋����v"�>��P�v�GN��dq�6� �5xCr�7T�,k�HD�b����3������I�^k�����DztA��.���C��^>��V����:�(&�f��o��q��{��A���g�a�/M9K���|�"Y�#"���`�� �����Ozy�GZ�޿=!�����)|�X�1��2<
�_۪�EV�<s�������i#�� R����t�|��0o���s�0#�=�b
�{��E�s��6f�aa�9��l�-���:U�1��,jZ�à��������뚍7d1?������^f�'��_�G�C�_}�.{�Н�_M#I�8����]q�ՓYI8�r	(�č#Bn�*Eq�s�Zhn&���њE��-��t˕�D���e���vv�Nyh�?U������Sd���[;cΉν�zI�>~;I��M֛f����V?�'��Ui��7=�&��V��3d�N���]W�?��� Fǎ����Ѱ��Owc
���0�_j�?]%��b��2�ц��(-+�Mb���m���m������zH��ӓ�X6t�~rA���*���5�����LLĥ�_��}E#S���Q�l���`��8bS�H;`�j�[A<e�ZsP��8�W� <M�s�-�^�r�7;?�k,�A�pp����.F��R&��H[Ӭ�vk:n�Ʉ�}1��G�v=D�*�]��)G�Kn���(&>7��o�2A����'����CpXn~V�q{Wf#HX	ޡ����K.6+	�P�X��Jeބ�K�a.PZ�$�܂/ki��AIa��&�ݣ�!��4�[\M���%�;'�����3��4���C�dpw���·�����]u�=��W��Æ�#��A�>sq~�5��o�+��j�xkL�cA�a词�4��A�Y����:�3l(2E��@���{"J�#Ah�i�:0�S?��H���� L!Y��:�F�U|��pG���Va�eJQ�'7��7�������7Z��S�e)�_Ң����f��Y/,�Dѻ�I�V�=~�%TɸV	�������3����R���C�[��"$�ٌ6�v�X�@��ݟ�ek�##�gZ��.���q�5������ ���*���_�)�>Yǐ��C�.�#m��n��!"�9���ə�fA�������e�#�Kz�K��N S�0�XD�U�#���Q߆�UT>}�m��*��t��q3ej��K^d��IM>��Z�b�z|�h{��:"칡�u?�p�x�G&���}�k�G�{�v�!eE`
dJLȎ1�g�RT̀Z�,��)3�3*h�Ei��u=�=�M�~o�;̮�V̇�X��-�P=n�"j�d���n�G�i*�σ��;W
eeU�������Tg��K���YF#~����Cb�ŷ�@�!�FC��o��d�?\'M��ۉ�;N�!r�&!���&�<Z�v���B}�#
�9��@�H��\��ձ@�S��WRD���<���]�����K쓾�X��KԌ���3��k��n:���S1��O?�����s���3����F���5&QU�=���l�O�(Ȏe,Fm�ҡT�c����^�c��i(��6P��`<�P:�����( cĴ4�*�ʓ�灨X\��̑�{�Ҳ�'W��$&����:Fk������D"���Tۼ�w�Hr��Y���Sf����
d����}sbB+HT���*8ʩ����{�Z���U� ���wŗ���I]�p]��+������d�4������XQd~��:@�K˩m��?�8�%j3����þ���uB�V����g�}���37m��'�4{hD��/���ξ��'%GF]�������O����G�hH�v[���G������ea�b���tCR���:�N���)��_�L@S�H��y��Ǐ+>�P޻�(_0������w�u����娴���q�1��Y��@�3�²�A�V�C�7/�X=��c?���D�.T~wF�$K�Z�w#���x��t=���`�G�h�k�#�i������ 6w:\N����w�)!X�^��
p�	�M���I��eڎ��{��p9IMg���֬A��@c���k�=[h|޾^�4��8�Y�#q�9.��
�%��!�1�V��������M���b�ߛ
n����U�Uydw�u�� ��ʷ��t���;ΉJ�m"�M6��i�G�����FW>�w~�c����ϰ얊���<���is�h�P�Ǥ��9�ٽ�����E�� L�4.�en
�ԧ�7�������
d��>)p\x�k�6�B�=u-�Y:�-�Ur���yW���̬>oϥ�BV���*DE��zy��B�
�Di]��U �`���%o�Fg�L���kL)%Li�����������2�����>E��A�bT&�Z��KA��%�Bwd�r_e<%j$ƀ+����ί�h>�=ّH?g�o���Yˍ�_��[����x�!���e��R?��h�E{9��.�P��jY̥��.��-���n�r�I栊R���Pk(9F�w|��-@h��Gb����|8�{=��Ю#�b���ڼc�#%]��))�� ��Qp,�K��m^<au������[�C�_G�����jr��zm5�����l������X�f�ey�>F�GRMj$�n|�q�H�B�m^����S����ju^��`$2j�[U��Y�~���v�����zB$�"|$+���� "�{���FCA���#��l�����,܎��X�l�6%�y�7��3\lܩ�~�)���G+�-�x�;���g^
�A�-�h!�F��[��0'��/��覽��,���Q/�T�w����ug��<X�󎼲Fe����]Mtd"AE��>8l���[��-�+)�h�]S[r� &T\��u�,��L�Iw'�ʲ���#f����O�P5ٮ�2G���3���C�,2��j���J�����n c^4�o�ї��d��e� �|KIֽp}e�gX�K�L�״N<D�
;�h0�zc��l�H��2��QpԾ�0��|g��}oN-��+\���}?�qQ������(cBBU�?6���n��8m>y�}��&�������C%�.o�Za�Q,��o\��-�e��Ә*���t.��͡RJ6���DEjL�KS��+���5s��.V�'��P��_���|[���<>�F�?��.�	������[��g��t�%�z�>vK#�8��}>l+�2>�	J��S�kP���F�G�kˍى�\؄�	m�;&{l1���o���^M
78_6g�Z���z~ �;����֥����f���kF�O�FZ	G�!H�m�@&�)����cN��Z"�4�^��05�q�����2b�����翲/�`����޸/P���ǻ?b��̚��:6/����N���^Q9�S�Ch_�<v��ID�t����w�x��JK��)N+�9 Yr���B��o;!DHb	�����r�=F̂c�,ʆ�T��7�%^HpphM<�����Cm@D��8���.�?4�q��ff/�m��ib��Sc�'ڒ|�
��Qew���xj /o[�/�A�>����S��m��R��.�xx�a�#Z!Nn�!�N�58���6�lU%����C0��-���X���%I84.�LY�v\ޞnѩ�;X� ��.��h�
���u�B�ڦ�;���<b7RM:���Ȭ�+o���t�`Yr�U��3y=�{�������S�!v6�N<��_X�����j��,l2D����X�5#�Ȭrz�w}#x@�;'�k���#�7�/>������G�����\3�n�fy���b��.�i)� ߐ[� O��/��ꚗy����e5�uU��Y�Z�Z�.��U)�@4e�eA���LT���!�[���<��v�	f���B֨�`R���F�;�D+b��f�nD������Ğl>oV�������L�&�/�����v��86׭&AL�b� �asdb�L,uɲ�4�z��8*GH/���f.���n�T>��DN:��$���uV�V��W�$K@�� ��<d^G׈6��3�x&(�X:a9��ܒ�t�������Z����*Pޝ������n�;u!x��9~�d/s]���O���E�5�c[�{��A엔O��h��V���ׄ[�l�Qܕ�id
ޥ/l�H���2~��f�H�<g�b�< -
�!h�rO(0.�+cP�(\�ź�w�i���[�����6/J{H{�dk�4�j�܋ۯ�<j���X�<��������k�D��%
�1s�p�L:��YN-!7s�+�o�hiÁ�J+ ��<d�)����ްI6�q�Η	�����?�lg�d��Z�Y�7�E~̝n�߸��kXm}e1�i��K�'�m��|�n�N0���ݮ��\O�帖�Hn�~��\�A_�&�+��N�����!h\��%���Gg�T�l��jx�7=�e��a���@�jdI��j�pD+��Q(�%	E��#u춣 �
�H�H�Cn&����TM8�H���c��-?@�e�{mٍ=��p»Z�Ɣe�B�Mb}!�����c-�>��%؞	:y.�l�u�U��}�a�Z;H��c:�&/�*��;�S�/!���`�NAifb�,,6]�"hq/p���� �L�A��Xÿd���}ƕ,A�%n7C�*$������I�<���͡eTޭ�Z!�t#���y:�ƞ�y���FZ8;~�q�h#�:�\�FE����<���:5Z%�RIO��܁%�sWK��.��]]ś\��Y���\k���z�:,�U#�N{��!E5	�.14� a���p�Yi���|I��lx�m��6�� R�����]�`'3+��侷�����y�����UN�`[)K�Arnl��,I6��d�mq����KN�☠�����y�3>m϶N�;J�7�	b1��pv�|K#t/��4|�`��#���}RG�94j�boO��LM]@`�Hrw�{��%?�����J����!��K��uJ���[���*iL�7�3�/�F�8�-Y�_sP��Y���KӴb�3a���=�<;��Q&r����䩳�5d�&�����#j��c��8	�72��˭�=��]^?�ݎGԳ�;%ѽ��bh���8u��E��!��}Ys
�8_�3ٓ���h��#F��N�+���"�'�6���h�K��k3����(�8��T�)&�y7J
�Ilx�ԶR�5Gu1��e���~ɭ��$
}�÷(�)2f�`Y�٫E��#4�}C�u�K�KD�Ma�O���ְ,�<�K�:Y�l�m�$�6"��0#�N�"�'I@�j���U26hZ��'�}CSt�1�1�nR�;��3��/����J��/ى|�[�?q�$Կ�2�U����i�J�3D����r��r޻̶�>i$�0%����j;6�$���I���K�����ތ��G>~�;�o� ���M�
��qw��m껼�L�X}g�e�p����6(Z��U��BGS(�,��8��R{�L{Y�?�|9�ҧY7��U�X�4ɠ�$�f���p&���o��!g��Lͼ�_7I�b`<7�C��~�N;��t^�7�4I(���\�T��\!�4���G&�K�&�#,k	v\��s����FNm��8QƧp/��+�A� �1���ƹ�~wa�v�2"���`���6z��c�6<�*O� �[��p��i���Za��.��Гߘ������� 	a-����]-�gh�7�]V�7Q���/��u����ysO8�\��-���n�$oeBe%�B5ͤ�zXLe־�s�M2�	�x8�^������v�{l&v�X9Rs��L���r�f#�Uv��ʸ����ߚ׭��h�3���u���<{\ᘩ�	W>����]��X\�
A<�-�Xam���*9a�*�C_o@#��6Ω-����(��I��	�a�9�����w�����=-`竨'݋;fS��oak}/�'{@>�'|u/����ɑ:���9,X���5�^rrp���K�~��%�#���-���7�E��7{Z�uH�Uj�=����f��X�05=����]}�>�P�{�D�7K��E�pQIW�F�Ϋ�zh�d�'���Ϯ|��&�����v�$/$2�f��ܼՁטq:L�9o�]�c(�1�E�gI��J�e�DB��#����\���)c��2���I2^��Y�-�=���O����g���ҞK�U&��箄�������bBO���^}��y5�M��eQ+4V�IO���^�/>oKc���%N[ˣ>�|�\���.�im�-�sNݬhy������`�K"-A���Z�2����_~^�E�w˽  "UbTb���c�E�]��z�S����H�A=��LSO��{�,˥;�#\Lk�D�z��=EE���"��x���6J�[�=���Pό�X ]n�3)�'���74�q����&RXp����=�G��AFK;�k;�8G#��w�^O�Y�-!�i;�G�4Y���⤉[�?w }i��T%Y7�]�RY�	yǾ�M��X:R6>��e�Ug���W���m��Ze�!mԙ�&@�o��*;�JC_����x��ն(�wƲ~d�I!�� 4�[SO�J؂�8}F)�}
(f vq����|Wi�����e�umEbИ���\z�iȸ�9�m4�V3�0���R32�^E��הK�����5�p'}��A#�
�R�zD��Ŵ�b`X����
��)Qi�#���q˅F9(:��<�ERLXQ9c{=%���@�#���S��!��g���>~�+%�mB�.1%=�������M�X6�"X?��4ظ}�Y8H#���g��Vr��u��ॅ��H��8iS�Z!�`}K|��������)Kww���!Ο��)bu��93�	��^�=28��f����
g�,�7� oI���ة��8%;���R:������� ���g��G�7?�^�L�,gG�֏\��T�հv�=uN"ZB�������".�*O>'�c�9�8�z��g�jN� 3	ALdZ�om�K���zNr�Z�i�Y��|�w+��T�����&�+��V�(�OJ3���am��1���)K�o�Z����[}Zz�z�������gw���@m�_�
%�K[+��q�s�� ��:��|K�$�'�9Wx�4�������Ӊ[ܴɠsU��T��v���516"SƯ��(�C��B�x���t�R�T��o��cB�N�۠���)�7�J4���h�K��&����J�TvR�(<��v�5�᭢e9N��%�tX���e�G�}�����u���?�c>�������sn��
��1�^��6_ށ�ǈ�@�%�l(�c�p�bk�7��/emx���[M �=�����#���ȲcZ����.��İ��3�v���W��r0k��C�J�����n�:��_�"�>>���+Ү1P���P�{���
�^�5���ܘ�����e��*��}X�N��<����{����+�y��h�x���+K�O]t�.���E��w��[	:9\n�����)a�����[�#4/���j�kh�c��b�1+�s/�6Ú���߭,3�~��χ����9
;��F���)��Q�u �A?Ty���T�c��w˭��b��D��vX�3�|X!�[2�t��'����d�@�3��%�QD�uM��V�e�h�7π���j	�1�Êm��_ � ?����F3R�O����3W@�Ep9��Ca%w�{�p8a_5	�Ѝ�e
?�v�W�,!Y(���_�'V�Qd2\${�d.K�q~��yQ4/�]���Zs�4���[���3t�}�Lu
Y.�m|�_<Ny�p�&���9���s�Ȟ�;H?S���HB��_��l��� ujz�ƾeT�6^��ܷ�	橿wdg���^9����6�M�f"�EիJ�q'��}vaY��P���X��)�M���Q�["ݡ��e�F{}����F"���ȴ���:		�(�cZz=I)�d t��X��?�ʼQL��D?�ylQ�fQ�{\G�)��c~�:: �	�K��V;�ȏ���\	����ѧ~>��E��5ߋ2�>��𢲻�p��V��:������3�~�����f��#L1h�&��Ȭ�����?Xh�5�xt�]%0�tIP9�մy��o[�mV!j��ȟ�U)�M�g�f T����X:�����-F+�G�m�ͧK[��6B�~D����x�|����;��0N��t���湱��Ǝ��=(NVnz܆�����y;�����a	�|>�1̸���,�)u���TU0���ɏ���N�����]О2�su��-�G����v}X�{�Kޢ��w7'��p��]>l��\��C�4��p�z�V��h!�.Y�ǝȣ����[쏅��cXK�7�P���H�}]fA���d>M�'�΃��֤C��8l��&�Ӫ[%��>#zx��u��8���h� .~��8|���1:=)�+�����9}�C��]�v�JW÷�KY0l���>��A�AX\�����{�d���}���Q�r���?���T*����(��A���K]��*Zr�yW���/xza�S��H���VM�o�����U�Z՜%�8�9O2�Q�����U!xy�D$����suNk\6��IJs�����Q��lK�G�b"�_���B��YiU �=��S�䮼��=Zʻ�"a���oA� )B]�a�.�
_u���_ڊ
����X���ۺg���{c=H?M�/a
ML����G����p��݇U�R$4�3�,S5�*B���'��)����
�/�pd|j�4�A�#8�.|X�2��O�Ʊ�K�NK�_�_s�o������&"���U+�.��|�Ge5v��w���w@��7�K+=�$��̕���
Gp�	!`�E���ǥ5م8��fD,-8,G��DC@m��D�/L?�Lع+T�#��U�1���d���6������{k'�~&"�6�=vC��ٹL��"vq�9۟rׄ��&�|�),h�e�2L�6LW��gU�dǶ%�4J5�2Q��(:N�c)�f�W���|���'�O�&ߦ]bJ�=1&�Pۤ�h�����g��h݆k&�G�/vb�ڜvEi���(o���)�9;ݻ��AM��OE�E�.|�%u��� �ҥ852��ж×bh�����A�����%*7�T}�K��]4��?+��X��}���D���Z�B����c�g���M�R�s����	w�pr����ݴhֹ�?��j�]��o����w� ��L�o��蘑e���/9L�5��V� ݝP2���F�	X���M�����<p�Α��V��d�6KJ&��*�ڲ�`��eqW( n3k�q��,�}�{�O�L}H����ׇ�<~�R��1,+�R�;&f���h^��ߚ�m�M��ڎ]�p`����j�oo���z ߹�G���F�:li1)�v}��/���8����	K�B�������bɘ9���{��6Po�I�jh^��إ(O��g���`}���J�T�b-m�xS/�p*:J�s���_񫦂jqZq㊻���QzKv� ����t����+�kO�"�D����^@������e1%���s���ݶ.C��>�0V�o��?�8rȢVC��Ա���94�6�n�n�[�y�,�S��A/B�����֨2[�Ɓ�$#P�����,K��V_FB�B� G�G�j5K[9��\	X�X���Ŗ�^�P���p����
J�*9�榿�\s-
n����r7� �͠�����t��!�÷l�}u{��"��G��*�F2X}�}��s�g�E��_�"ujh�W�V4f��<Wg䥶���.������a�Ŷ�ñ(��]�0o�1<]�n��b�ɛ4�7���+ �T{4Dh�3�m��h>���;��Sc�H��~�`��%#-��Z����������Z$b������ͮ�L�$�/� <�^<�[ۙ ��/V�W�Zvw�w/��׵T����a:�2�G�P�1}��V���yb���~��?�t��[.yO���g�y=�"��4��Pަi�S=%��(���V/�~�%��/Cv*��#p�6��p�k�����M��޼�㤫#�,��\��	bozx��`�ո��o"�C�I�ߛ��TM����5��j?�D"z����z�ơHN� 6ҕM�Ɣ=Q���~ra	3�֦�N����W&���6Y���̓\����[���4�Dߗ �!*s�a)�s�cD�d�s���ո�� �@�5*ʃ>�{ƕ�B�ڥT��q�oѵd6pf�*���s��N_Ew��eB�f��~YԨ�B���}uu@x�`��zq�A�U�����I��,��������&�|�V��5Ą�e���F�����G������ի��Qgt����[2�C�m���ݖ%��
���a�M�6_��d)�'Ä3焵��O����[�od��-�\R�(S�}�����kS2���	�p�8:�[w�[��\I�c��r�I��>�e��eT4�g(�]*��݁�A�*���7~�&��M]"=1��"m�ط��5�V2Pa{O�6��V`W�q2xӀYI���i=�L��eג��sژϷ�qj`ͯ�a�3���æӜ�FW4]�E�+��,@�b0Z��"��knԈEՕU(o���m�_&�K��M�ki�����X�[�6e��ӕ�]�{�|9,Ȣ�s��gw�b�O#s�Η!��+�6�V��4������]�$\����DIX�~�o�:(D�:�e���J��Z��q�i�|:�a�>�!�fK�4���*�<���0�-L@P 5�ҝw;R~z�U���e����`��[l�)8.�$� �r����ԋ����<��^�e�n�u���O٤b�&�oɣ�d	K>C钙a�r��F��}F����Jm�����^A�� �yCk�
��U*h^v�G��_3#��)%⧌@lT$l�ߍ�t �&d�ک�G�:`i��A��c�o8_�;i��OQfq����Dl�g�L�Y������#�\��m����5d�t��]ǮSm��|:&�'?��U|�$��3��L�^���환�B�K�b�	�8�g0�N\���Z�t�S�BB�h���̞��1�M���p{�Q�	�"��s���Y��Cz;Q��2|��EP�gB��FW�a�&B	�Ȁ�bd�ˁyS�<�pvp�K�h5�ź������,�����cr�?�G��%_���Vo���+�380����A:Ș�V��;��*�\�E���s`��[6��}|��T��&b���`��A Bx5������c�E�o�m4�i���$��⑚����%��ᐠ���l����������'R���Дs����b� �I���f!.У��"�%����SBi���A���Y[5�Yv��O����u{R��q�߹P�&]�$�W�?%�?W�%�m�*�B����c'%q��tMqw��?���$����K��B��< �1p���J�1��xb�-5�ĤͰN& ������G�k�.q���ye�a:%�Ʋk���$�mMe��u���Ũ{�|(�����xŬ�]�b(Ŧ]�Y�	F�	7��#�P��Ԭ*��l�vSS����s'?�&��>��Bs���1����r�;�X��{�b�>�J�pr��r%g/~�ڬeE����>5�mb��T;��Z�E�}��CC8�ٴK�/!�����9$	�J�x��bg�5lo�>Ծ?b����~�͖5��+��Q[��Vi���q�:h�ȉ%}�T���kk�Bo�_o	�ΰ|�4��8A�_ �W�����{�?Q���܌Q���A���N�C)b�$�ո��p�_Q��ƞ��[��x��ڳ?+nx���f|�q�_?��Z��v�rܥC����j*b����v���m�9f<��.�;0�xǨ_|~!N������+�ŏpN����X�k|�WJ?�h뭏U�O��|���d�|�%JF�k�3�n�/�ޤr�N�6��v�s y�-�
&`Ż�s\K�C�+ͺՃ̝�[�!��d{�zS�V�¿H��\}tF{�˘Y���Z�!U�_��{ʵ^�r|�ԏdNS���ٛM���߅�d��e��j�/�?%�D0I렽|�Y�t�%Tr���}��j��OE��be��Q��;��A�&s�@�z#�^0��Q�R;O�%�N!�l���ӒV�HM��HԿ�ژh��^�K<��.���+�[e�W;-�a:�d
`��0.:O�E���&~��]�U�,;���.|�.;xxe�-Y��/v7���M�9���q��Q�D`�,� W�ul�e� v���O��3Ƒ��|8���e�Җ7�:v��|n�t��SsPw}��|-��/_e��~��|�����sܜtg��4��M���6h���WB�?2x�}�Vu�Ӌ<�׽C���� _	�<�O_��[!�4���yK4 ڸ�z�:Z�e	�H0��~[XK�9ZS(�	�4�F�U�%K&jڴf��`&�ɷ�۔��$<S;s��4��Q� (��Ds�0�o�l?2Q��j�U����tK�5\������=\�m(�[��ه�\�����tB?Kyg�
F�~��~�s����"�kYT���U��՞Rs+�;5�6�*���F��!{i�� ��Y�S�N�����������E	�Xp�����-?���\!}b� ����DŪ�=׵W�����尤�����׮�G7�4ʖ7�!'���yE� ,�}��&�܅k�?��J����4:��܏�e /���U�<�12!T�	�6���*t;�#��].6k����Y���fw�M���b�z�f�[������6;W�,��t��ޜR�,7�&�!Ƈi1�Ȉ�O��|*�рio*1� ��U��W�w���+Y����C�W�x�g�T�:���[R>��SU=�Ъ�=zR�8��ɃhK�a,蔱�*Χ9�[;���c�ø�_`�l��Fn=�;��+D�M�]x���@�3���0-G� ��4�P܂�e̷��L�I�A�N[	!l��؛�!���"q�OB��a<A-�_�8���p��ˁ>e"�q�N�MX1ᔜwy��iq����	5��	�,�$_�2���1	eܑ����ex�����W����F!�Yw�5y���Te�L3�k�>E�����~���m\6�q"�х�`���㤓�.���U!]Y�ɫ����w�8lm-֝G�lDƃ�0;��f6��O�����3���T笽ETW~��
˞��C77v�1"� ߗ��A�"���S݃u$P�5��3b�����Q�g+��������@��Y�2�d��#�:S,-�HnA�
F!,޻��R+%�f�~�;ڣ���]��KK}�K��~�U!,�B���r,�Z��hr�7�V#�u��6he��F��[Ea�{�U�����`耜GِVٚ��hu�Ɗy"��H��-��}�X���%��+R?�wd2˩N�����s/���U���Xw�q�Rlh��4��k��a�E
�����ZE�MȜ쨸,�ܟ�b��׳6J�0���2�NAL�!���`t��!�)I����b�Vm%�} Q�'�-�n�Rp���][��Cl	ɳ�
��:>S7�����`�5t�I�G��{�n�(�uH�]��wPr�̡�bB%���\�Pm�"O2��OR)�i��,��"`Kk�&�4	S��K�X���n|�>c�����Di�T�ժ�Ż���	cXѮ���h�1'$�������\���m��^����?:�+�#j毡�qeQ��L+5<Q8 !��p�_�*5a_�E���x�������-3��p�f���j���aBxk��ëi̬�s ,+C��21co�������Yh_�������t���]�`�����f����/�3�z�ĩ<�%X�)��F ��قh�i���PՕ�S�P+ ����֮2/��W��M��P�>S[�iĝ̣��=F?6^zd�-�8Z�8T�W�vN:�"of\���phl�:�a���}91M���"?�73o]�mT��_��o�І��c�(����%s�32�����!`�7+�� �I�M���?��t��؊~��b꽔��Q�F�~�eTH�ж���S������)
��)�ojJ����[Dr��w��	�k�m��!�3A�Di�O��.��WDd���+�B��2�
Z�C	[l�eP�VORk�l=���6q�۸S�X'QMBL]������^��7#S����r~Y��!j\eq*vY,��GOoy�}�V�7��5v���E1p�� U���+�3�Ϳ@5�;L�}�z�'b��+���_{�`���>	D�ɞl\��+W���"���C+nT�_�>����Wr�4AAF�$�W4G�ej���{��(:�K�)��^>��}���j��о�1j?7����I��ۉ��E�� Gkן�H��X�m}/8(�5�0�B�߂�B��Ԫ�R#�>(-U��&�7���X���K��_4��-t<s�iB��\o�À�Z"�2�I�K�%���J��U�����ky ��=��Gҕ�ԝk=�|�ӛ���`����"���eJC�t�%X���\ӯ�Un�(��n�.u{�ઐ�wS.f���;@�9��~n:����UR���d��f�M0Z��^?�FX��j�x���d>c�Kw5��Y�tEk?~�j�g�+aǧF��ju��k�W��p �pL9�ŉ3�Ƃ�f�MW߻Fa�'��T�/χ\/����.6d��K����C���������'�p�=�'5u���sB�"*�Zx"t��l���$>�xzA�o�'A�s=�G/�;P���eɰC�B,%�0��8�+��LQԊ�98l��\�l���5+ ��i����e�+�	�7�x��IE�f�
6�!ċ弹Z���P�����M�78�=���h=g�����7�-��~���	bBm����iܱ�jE��>ׄ��i+cMf]WH�tG-e��W^1�fnze\ �?vp��iO����**��"(� ��@n�;hWV�Z�յRx�f��/,���7�aּ��ok�_��2�Q�+Z��jYŰ �h#F�(���0���C�`g"2��ސ���XV�ro��Y���M�,$���{Q�{N&�7���N������'e|�@CP9�T`����%��5�>j����Rw޹��5�c��Ts��Ί��͌'�_M�H �#�Vɠ4'�j�z����2N��S] �t`��I$,�؊AI����_�xVGw�������	N�;y�<�yU-�D�zy�#����=?`0 }�t���?����)2|J��:%1̪���V�Ӟ@�e��WC�������3W=y��	<�ɯ&�JϜS���S���ha^���_�D���ل����45���Di�Q����/2�}+6a�0�f����~��6l�H8#�wε9�+�T���~�y�h�s�a�ܰ9u��:�����rG	3JM�]ռ[,�D+r�}+v5_���>����q���3�Z:):+���~�K��\ȃ?��_�Q;O��'�:�F�]�J�#���m�7@x�"ET\a�P�,*�L�-}������]81�<V�����d��a0[6K���?���m�n�>}�0���N�I�-�I��Mo~�O��S�l�2~O�Mtt��|aH���d���n��������>��O_�d��Jm	s6.�����M�z3��5�d1����1E=?_�V=Z�g��4�e/��1�� &����Z�U��Dz>����@�����|�3MӬug�OƬ_��� `����h�PB�s+.�Q�R;��?`4_�@�')	����S[ȵ��ja$ G���5����YH�	r`�۩��#���ŗ<$��#b�{���B|e@��i��u�U]�j�R�C����}ejp@��j��i�p?t�q'FXF�~��y��8(C���v�{���b��7�z��ۄ/EB\��.��[�c�򀜫%Yy��	��ԝ�x�2�)%�S^�@��̎QN��a�e��r�aݭ^J�͇���<�s��^=�t���A3�'#m��4:xg�u��q�.}��d|TY+�r�Q�6Ƅ{.5lg�I��
���_q��m]��]ؕ1���¶&�(�zm�%n�h��ؗ>r��p��l5�6�Z�B��k�	����2]�#�ݨ�*����*�����ŉ	�'ԢY�������8���z�R7�Z����iJ�	�Ma[y�g�����ך�����e�ԢvŨ������dsZ飝~��Ί�*�e(��o{�.��6f6N���[�!A�z��Z��M��1?dm��S�6�O�~��Qt��ZO�R.GBU9<�c	�nC�m�*�睟�~ӳ�/�=l�um5|�}��<E`�n^�T��a�y*0cUg ��죲��r+͸�,��Hɖ�l� �������P�=;�l���Mxo�Yٓ��egN3����O��>�g���ء��ﺰݳQ�OK��$y��(CE�nmR=#]2#^��[!݂�o��<����JȈ�LzV��5�c��s�� z�k��m�x~=/��x�-8��e�4��v�a��k>���|�a��*�"�����J*�O ��(�R/@\������������!����D1d�O+%���䶯ψt)ٖY��I�u�vvڔ��q�mW~�lLA����P�\�
�O���i�p�X��t���P����yD���i$]�g͔7�2;H��y8r�S�v��@	M���G?��Y�Z����8̗m�4������Q�Q�����"�v9���F�M^�;c����
 �	�qZ�'rr߰Y�9����M#Ja�~+}��Fm��ܿ�m[z>�zi�*���&;>HS�e��L�U`)L�k����L�ߚ:��3]7c�G�[�q%���ʨ^F��<s�8}8g,/;�� A;�z�X�'����#[4��B�C����'����aT�=:��k�#j�a��׭�����7�_KtuX�Ϡ���T7���W�q�� ����-V,����(	�*�F��t���w�f�� 8_Z� 7��4�-�x�ַ��}��f{�1���+�0n��f�q�^��)��B]���J#���A/�v��O�Ӊ�n;�	�IYkO��&<�f�q�I�p��y���s��T8T����%]����;�����UD�>�%����$���n�C�SP�NA��A�;�k���~o��?�r�yf��9����h8�`���U�Fg:��U�)'�_?���B��E��$�����nQ�Č�V��Et:�fa��{j��k�2���u��S@v~|�9���vZz��9<s̪I�������u%󃥐��CʩԎ�=&�@�[󠊂7�O}�� ��
�\z���hU�̝a�Tb1�)��}�4�Zl��$��Ky!��vq/,��Y>Hv�9�)ZπzX�C���B�M��u���c�@(�M�)���s-9m��q�V�H~׾�7��(��k`���Ic͇���`�T���kM�beP�@M�yH�V�&~.�����q(P0V��%*�1=';�y�p��%�d�U5�	�C?�W�3��6��7�.��؜�F��l�QR�T�Jag;Zӆ������|_SkǅS���JBV%�K����"WL{���������3%��|��.�v��,֤���Rg��S��	�yVc��P��Ƨ�WRe%O���Ԫ�7B��Q������5Y�����2ʞ�^a]�n_)%a����ɤv��I��5����m��j�YwS�@���n#�l���Â���`�6Jq�~cѨ��ȝo����,J��a`��'[[ķs����)���Fl�j2C�mתו���L���J<g&���g(�X���Ϯ��^�]۝�5��^`���$7���,f呔w�F��0KvE���X����ͦ� �ke4��n��'�{����ۄ���ӎ�-dᖸ5c�:��|�,���w���k����U��m?��V��K��(��zx��?A{vt�3�%}Ѥ�3W\�l�����M9���ٝFX䨗����2>�L}	���u�c���c���T�FO�����[+�&\ � ��>@{�"���y$�	���)Ž�����G9�1x�=.޵�9���	<�vo�U}��9/S�����i�!�yHYM糾Ox5�A
A��E����x#�oM�Eb���uL�wj���笠4^?�Q���eT|�A�G���:�ޫҒH.��~4̏k?%m���u�U:�u`���H뫣3��ͯ�Z�Oo?�>_T�y?#taT�e�D��od79@�AU�v���\}�EK%�n&ڎ��K�2��;vm��g���A�n�#���A4^\Dhx�R��Ւ���g��Km��Q�΄�^��y�x���V����$j�\��.�ћ��G��2_4UVd�54w+>��W�Nv�_����<6��������7d�ٝ ����b5���\J��z��Po�9F.���V�P"s���x|㩟���Քg�ri��)�B�^O�g�_����#y��ۖoЕ)�h��}�J�)c�Db��b���t�hU/��OnfsC#�ZjZ��;��̦.��>/�U�D��8�F��U" j�3Y7m�1o^=J��ׯ�xs�L�D���"�!3|˷z�NjѺ?C�p���ZZ;�~�[��"r<���*|+#Nx˄�L�O��u����LPѢ���v|��?{2Df���2- m�G�\DQ��ok`ա�ʯ�Dc�Z|ь�^#�m>u|���Gb��q�_��|$ꩅ>XK{�I��㵣�$�/6�$ۖ��0�K=I��q3Z�g��2A��J����Sg�|�w��IT�A䈐� ��w�]����c��űO�?`�z`64��sVE)>Cʭb���a�ԟG�>�|�h���5�N�vLu�o��i�~yR��bDN^l^vmD��F}@�+�Z�x���I�@ԙ��� ���a�zb��Py|����Z�x@���[�wO����H8�e�^b]��b(��5"�R��]ux|{v�&?J�������^G���_Ӏ�F�q����vP�r|ٴ哀l	D��6��
0��b9��3ͱo�b��P��04^�h����P�����_i�"
��aH�:���~�)�4� �d�C�t8R��<�f�#�q@J�0�{�����
,��Uj�����Xph~
�^2��S��2�o)�ѩ�{2�!��D������>eYXğ�>�D�>,h�̂~A��V#dq�Mh�hK@B�w���v摒|:_��5CE��>�m;�M#�3K�U��AܞR@����B?�����+�(��
��笊��4V��G����DɄO�����OʯVˁ�LH������kZ�עmِ{q|V�<�R�%�%Ҷ@[�+�����M�H�(;���wGZN?�D�l��
�z��$�7czEyw:wl+�/�������m��#�_�g�a��9��]���@ꨌ?̭�"	q��
:j�h-C�DE��� u|�Z(,7|X����T��&�����������y�i6��ޖ�]��|WY�,�^�N�
�s)��`��xT�(�"��k��L��R`m�;M}٩����G%c+K���Tz����,��X������ǎ�i���]gMTYt�5��Q6�J�/�Z�t{ʰ��7��e�j����E�P��y�S-�ܧ�Ʀ�����Bi����
�׍6���V�m� �:�[H�d�1��6�D}ѐ��gA�O�ړ�Z�JF�?@��	�E&��4y�9R0�(��&�M#^fgX�5��!s
\�?�L�����ߍ1g)H���3�L��F����R�m�_LM��#\ O)�ڄ����mWVp+`�ߐvn�*UO��L��gD�X$!�õ�G�j��c�i��9]4O7i8�/��5M�]� &�Y����*��z�'��W�l^���I{�0�E�t���2%Ҷ{�b�f��G���r�
��\e�B�%~���Z�ax�Rg���&u`�|���%���~��x4H;�g���vB�C�UT�ج,�._#z>�*�m�/0=���QY��&#n�F5���`��}$t�s���7��F��e�b�TקB8(��Fg��@�(�)8�4-��
%;����ˌ�?7]H��@+���,���Cpwv�����m�В7.*�y��q�6��ؔ�藉�J�p��M�V�)x�n`�F�IZ'�]�?/�	�V1ԝC�� ݧ�F|�B���F����[A�l47�˽&���w�Sc�[��Smx���<��\�uJ��9���t�y�2����#�[wP)A����N��)���"���&.��#��iz���`�dv��%�'�ئ$��jC�cQ�f����l�m��(0�n�/7GS�K�d޵���0�F8EbP�����-�	��+?I�p7�@�fO����d�5K��ð`��v�D�cK��<fVN,a��=#Q�����seN*����R5���@��L�N���'	l̋��g�V�JU��i�/[A�_��H�K�-�3ּ�Vq�!�h���C޷&�y�W��*	]������72'YG�+y6Y���*��"�W6~��7k�b�z�M7�(�a|�uv]z#����Ǚ`��f&�����`Xⴧh���R��.���ň
�s�:�.� �:��%��m5����۔�qk�ʒ(�%n��;ҷ�\�F:]�������jϠ�=*��[��A,�J��8�Ð��[���Hc_S9h'<�_�)Eӂc�02�ŏdR{�vW�a7=���� �~��!�e=T�	5��7����3�¿�����#&�|��W~�G
�ZӢ�h3��@�C�vJ]]���E�{�����y�LFM>	��y�N0��m�/�Ħ������rX�c�~	s~5�{L|u�P|P�C���z��o�D���Z�����<��2+ZK�h�0Ȟ�*��� ����g"ъ��bh�����AbYX�R�qJ�,mt�`9�f;��y���N��%!X��.cXq� ��\��'q!Ѐ�x6H*y9���#��%l�^o?�E��3�:l.�l�[�ȿ��V�*�h|y�����������[>���!���^�Nsz<����X���WK�nB�,%(}b�%~�K�!�95��.�{� ���}��prG^�e`t�6�˯�{,�r��?��q��^��,�8�t�ޑ���e�_���9�)�n�*�K�%�����+��ᐮt�ֵ�_Y����L}���8)Ǚ��FZ""���6=�m�
RK�ݍ#�̷��B`gAknZ��Ú$$5�m��Lhn�}X��`�e5����O-8�NOV�����×d�嬪��R��M��K���^�D����;Q�+̐����{��U���?�Ǒ�F6����8~'��N����q��^io�|��XG��kۆ!P�uP���n}���辺F���{��/=Y�j��(��r!3��o��ד�����<�K�9b\6�-����t�y��@FPlg�Cm%�#��OI���w$����qPh�JN:'���W����`Pi��܍3�Dj�g���{[��R�W��>�eqFɗ$R��\�5���,�z��>^�}�xSj)���ۃ�U')=6�"���RNa����#�B���4�Ugf	���H[)V^����-��n���r`�ltٲ�m��Y0nOr2C�n9���n��em-0.��V��kѼ��[Z�.� ��c��1�a�Vb��7ڗ�������KI�ks�iN�M�D�PR-���Е��Ȓ�F'PQ����"���S`��x��ZA������e繦t��d3��_�i� DHe,�Nss.�����b\�$�5�Ϯ���M�x,����29�T����y��ړ�ש����j��	�x���vg5?��{�nk�lb�EKߑ�̩�+�����,3��ZZ}��%d�פ���0&��L3��|,��ɳ��_	�}C���Shx ��'�솃����j��E(]jM6+{ٔ\uP����[,�֟��? v�-�ל�`��d�M��HUƤ�p6l :0�ْG��#�!ZhiV[�C�O�+�>�{}���zK��n7����>6�?M�U.r�Uj�/䌴�����U�b���J�F��v�C���!%8�<o$�:�E�3�9�vD�d�!X^4�_��΁J|�w&.U��Im�iz!?�\:E�&4�L,R��ǱG�0P��6sQi`���oӉ]���hHn�:S\f���a��K�v��n�d�5q�_lC>�(Xx��@T%(�����`�e&�CR˺l�6��g|�LnU��+��3v�J� �1B�o��Yn�6o+��^��0����ൊ�^ ���0��s	X�rC��;h��N��ԛ��X�Ds�8��#�pb���.���9��]I�Ȓ�u:0S�)|��O�	,/����1�E�,f����1���_m����$��t�=!��V� (�j�}KEb�I�@�P�^f4�IhӔ���gd�������|6�� ���&uH:a�~H3)B��b�v�ͨc�z��&B:��b�NkS�e�_�J�C��\�����V��"�=�a}2�q������T`��<d14�e6C=�C&�E=dG�j����}���4���Y޴�)���KjD`���Ĩ�*�;�tc4�(���;\T���НLE��'�
n��s����s#�d3 �������8�S�9|�F��'��%'@TA��x=�����10�'���6!8XF��j46�ݖ@��)մ���S��h��n86��Y �U��R�����a�����T��!���M���㇞�1�+:�P��쭱v�͋xؿP����(�����Y�0c��2�R�=W��i2�7��͗��L��:�P� |<W�w��l�9�Ζ��-��}u�93J�ߨ���>ni�����E�k�nY*8M������\D�S*�ҏ�wtdNl�r��e�BU�^�^�.�_���	|��{��o���R+�L�n}��:�5��;'_JuF��?>�Dz!�C�_���݉ף�5Kե�Uz������"�w��z��٘g��9�c�Е�h��7|'I��vs�e�����E-��/������E�J{�C���=�I|qua��i-�^1��pk��Ȏ�[TM����8��6f�~ʤ½bk��R]����ap-<�����vr9sh�*��Nm�:>�-	]#�!ȶ�)����*e�ǂ�n����F����E��ԡݸ�,ˢ��>댑��lQ��lo/���ԃ����	Ϋ���;F�'��m�.�
��f�?9��n��ꕴ*v��Gh����ޅ	dG�	��7�����K<���5����\d�e�g�փ/ّi��R<�Q2�-3P��6��8J�v�ֱz�N�A�k|�'E1Ւ�d�`׭��C4̆�ۭ��1�@�bI��;�n���C�4�s΢�s4�9��M۝Գf`N��t����i�_�o�:.�����f�2xܾ��E@kjehj��������dkO��>oFM��o��6��a~x�0��!0�[�6��{�K�����g��bF�=�n�	�l�nT���S+G"/�za����g����h�ů�>���B��O�=���(�B���G<;�(���"�y���N|Г���Hg�����w1{DS$���t-�8�Q+={ن�)Կ�tW*�)����ݡ�E¸=����}��p���
m�p�´�p&��?8j�+o��/`�ԛ��U0�|ZY�M7D9U0&=���a������k���Z΁6π�W\;*�ԉI2<��O����{�q��K"e�	G���AJ����(�@<Nf�&���'���+���]]�� ��Aٲ����KTp��<;8t��4&NZy�r���b���vY��ƺ��!b�Kv!途z��m��X��6�XP3t�=��`��v����q�j��¼�%��Pn>e��N�G8]�.��w�@U��ҍ�/e$��m�U�ފ�6j+P�n�65��74�%����}_�Dh[�ͧ���&�����E%��J-��j!^�rS�9ԙ�G+�k��5�KZ_3�6�횴�8�χ�,MV覒b$Q�4�9�Z�Vk:��=����%E�Ɓ%g�Mϖ�;��A{�4�����VY�ں�on�l�/��p|z����7��ٯ�6BV_v�c�	�Mc��W�"y}ţq��{�9�[�`�k��%R\!�Bw�A���W(����j��z*|]09Ф`��f>��ՁF	���n����y�=���t�W1�њqB��b'JHJP<3{�H@��^�)X1,��WU�߄>�u&1L�?���;R��ɨ8� ���qH�C����j ���=�M�=�(�5���*ͥ `nS|3��9�5B��0�`z�<���ON�f���@�y.���E�X	�U$�����&{=U������A#M������P��Iͩ:��Wa�6n�(������ht����4:�G3��UX�F"Z w��}4�~y#v3�k�����2��L������#����ԁV�+:���]d���k�L3^츚6i�j+�۴9J������n�I�>�%�.(6�1,M$���"1_j0�AiO�J���ґ�`�[���d#VLC�ݶ�cZ%������w�ƭ�fA�eW�As������[�2B���c�]��Z�6Z�Ғ�hJ�p[$S �p�BF𩸉.t��O1���*����=���4"y;�C�!)IfE�[_U6�)f�����[��F]v�����-U8�mp�ƼS�������~`�l����*-鳹.r��s��,`��$g{��Cj�NU8�>H����7� m�`!�i�*2'o#M�C=Ιg����Ǆ�3�ϗ��:n1=�|����a �~�v�����,X!/\ҥ��� ��[q�娽.�0EW�;G[-i�+8�-�kxQ}sJy@/	$!��ZYџS��nY}�!�U��d�w�Rlఋc���n���G$Z���{uoƹ������2S�J�E�g������D�MU��#��B�""����I ��c]�H�Rw�>��K6�Hd��
IRHi�b���i��藈ic_�Z������!�|3m��@G�1�D��05K;|�SO1��Ͽ?JF0"�����Wӱ}��'�a6ݐ`�T'��AiRnX)����B�L�B\�J�6���8�Rc�x�ˣ���+J��1'�̶t�(9�����<�}W:�t�,�Gbv��Ri�	V�x̵���`��E$����=Cd|	dS����B�w.�i�3����Ki"Eψ
5�¤R��<&����5��N1�����f���K�m[z����ry	�Y�ZsIdS��PxM��i^��|��]h1v��K��,v�א|t]	�3��|2��\2��DG1W�������_[��z��BB|j��3��]�� D1L�|Ɇf�q�W�h��a��E��2���D��ӈ$�6,��>C� ���a�|<�Bt�����4	&���Z'��.�zG;���V�pǶ��>��`M�������� ��1�9�����Ӈ��A�`��Y.+��х�t�2sb��Kn-(�w�|-N�����s-0�*R!�'f�"<�G#��D�-�]�&��	�!�$�a����k�j H�Cݵ��qY}�ƈp�w{����xI��ψ�>�یt��+8WTZ���^����H��]�����$����Za��GWWPȤ�2�����%=27{Qy�%�"�`�T�s�N�ϭ��٢k3�����I\KvG>��eպ�d�Q�^��D/�$��^�o�궋��*�^��wա���>[NC���e�����=�l.�K]5��T66�ݦ��e��ҽ~=D��&�M��Sb�����oę��y(�G>�*��<u��ӣƅ�E�Sˍ L�4�����Kh�o�������I$B1��וj\�>��Ǎ�!y�~X�6�m��~�xA^vZ��?`)�7�UY�H�-�:J�hg	뗄�"L�h�<8M-��P��;oٮ3)3�J���[��݀x,&����h���"tک��N���'�7a�;�p>�I6�x��Ƀ�VJ[5L�M���٢V.���}�\�cX����
$���}
@�=��am�/	���©Ce��%�J���F;�ǳČ�v���ܛJtř���Ȭ-!<y�|_-D�~���xA�4��h�n�:o�"�A+U�2_��>������忁�t������X��(gq�@�=n!���D�^�N��fIK����D�2�'sw�Y�t�U��5L�?x2�z�ɝ� 3\���[�����i#���=���0h���q��ߥ����O`B4H�8��_Y�������\݅NV��M��ػ:�A��R�`!92��ݠ���Mp�i�k���m��x-X^^~�g�;�'�;5��"i��9c�.�3���/��A?2�֙�ԒڄDS@����mQ�m�/�9t�J^Se��-|�?��_Ǉ*�{���0�v� Qtl8�.�ܡӼ�jF�5��5{�ܝ&f[֝�ҙm��K� ��~�h>�k9�	�XImo�s��w�^��5H���t���k^����D�6�wJ��� ���0F�mqX����!�\�8?;|D�����kL�y�d3�UYs[�YVy��v��5��W�F�4A;b����\W�ak���^H�pj :�12p�b�١�S�����d�jG�Ys��ϷG(��ڍL:�oo]��Y��c;�w�WP%�)�?K{�T}��������學0z=I�6��o�P��l+.��ɀdh�{���2�����=%A�"��%�
0������j&����r�ҩ�(���?�����n�J0�q��V-���-6Nӆ��^9��`�o���m�ZKM����I�a߭4�ϲ�+�f0d$�	W��SP�c�5:�c�0f$���,�k��Z�V\�y��읆p����W�����z��0cSB�k����xBB �����'����(�GMA~b ��g_�&[��8�������H���^TD��y�tS�Q�s,\�1�6�nQ�kg?f�qOѱ���-��F��
iR�Yg�"��%d��m��@t\�v�lnh {�y)+���E,���Z��;�~�w��M(գ�i��鲚��E�*鍂$�Π6��9����s����v屷r��1x�R�(�R���nZH
�^Z!x� �Z����W�('�/��r)[��n�ۄ,)����^y�j76��x�^}}_�_B�E��>}@�ب�f|,�	���_�ϰ�ۅG�#�6$�(�Ev�������Y�E�~�j�s�l��][Nv�n��G�/߫E\]�)y��~Q��d^智m�S[�U�o���������pW�WȺv��-v3� �XW��rzKdE�'��c-�HtH5�Hw.�/r� ���T�!n@7��ް�hs2)@��K��(��Pf����O��+4�;Qo
�(�G-�������nӚ��m�U~�>0*-¿������D�ym��ph[����M��󦹵 ��Lv�;8��p���۽������!o���f���ҫ���c\Z�A����h��
��_R*\;w�����;�/N�B�x��ri�4(O��^�W�g�-z�3�fH�X$�Eٌ��yg79s��ӱm�UM�Oc�6�Ɨw�,�]1bh`WR+�Ƙ��c�]��ο������d9��Qh�34��Ȟ�>���bC�=B�+�-�f(n�D��V���+m(3>� s�:��=�������:x }Ñ�I�}�W��/�/���_�����6V�ur�twJl��+�!bN`��M�c9m�dI[���}��_mQ���%Lǋ���~�_�4�:=�������Oo��p��V�+T`��S4��n4Þ��x��^9>Ǽ|4�*(�#\Gw���q^�"��9���M�8��6�����؉Ij !��ʌ���D�a]���!	�ر�J`0�ʖ�fˮn~C�P�j����Z���y��qA[��1}s�C�/?ǁ@��Ĩ|I�y҅_\7?a�CX��#S��m(��'
��y��~�?��8�h׋��0=H�f��@����1����Ex�J�>p��'v�n6���T�+��)wA톗�����������h��99�B�ԬW~/�:�e�G��i6Ue�<��U�6���'ڂ�j!��! "�W�D.�� b<��RY ���Elŗϛ�֟�T7,��LB��eN���r(��x_���Z�~-��%��Zw#�K�,�Zl$�i@ip|�e2��_��	��+���J뫉�*��K�Z���}:�E%Ǡ���=�9o��A���zۼ8F��o��%���N2�)�7˒�F��*�����|KAj�uV��`��n��!�O'|ٿ�^��V�n��+]f�n�n�~X����N^]� �}i$Pԫ
����B�6��PŴBzd���`�:�[H�/?� �poLP��B���E�m��|�ϼRT9E~�_�	��o<a�B��D�ԛ3��v)����ڵ��9nN�&�4�o�:��s���.�
H'KQ�-�y�?CNX�n�=Q�c.ȚK�8˴�y���*8b������j�ҷou3p���vN��
��6߾h�:�5��h�D�1�d6�C���$l׺)1ŸF��%�h0.>�
{��L6	���\��hr��B����13�ߢ�AI<�ұ����ϰ��2K������&��y��g|����ǥ�`�BFP?�C�u��AL"S7lp��B��m���mcJa{��ry?�)>��A�7Bf�M�����ODӮ��w�ڨ���B���7`ݘ4:I�l8#̐���5k���y�샅������"��$�PO�$� ����~Y��f!���cp�4ԋ{�*�������F�J�0dp#�pF�1/:�:�J-�z��%n�|�ի�-HXTa�K��g�_�]�x��e4�S0���5�����ˠW��:�����)1���_�]O��2	0Z�c!�;�Qq��)���9�l8Rk��|�-��>{�9깎4�^T�v֙�\�	����wmu>�y��c"��m������t�/h�{}]�Qx���)��G����H�@zU�n�u^����u(���[]Z����ɎǙ$d�Т��k�<��W)�����ܹ٣&2J���j������>�����7�:T�Js�C��C���5S�7��x@�U���R���7���^A�N��|������+'H[��S>$�'����s֋�d���-�1+�_P��~vk��&���soz���2Ρ����!sm�A���[�����w�����w��A���t�af-�E�O�l�}��Z�F�����M[��8m��J�"�܁��:�r؉j�'^��t-��R���`��'L�lk�:]��:�����4 ɩ$E�/��dZa�3/����'>�$��C�d_D�I���)>j���d�A���X�)rV�J�a�6���:I�����8��+�-X�r�9�I�qz�������a6�tDh�J#ab*2���2/�ٺ��5�nH��)%0��d�ĩ#�7`��AsT�q�b�G��u��3�3��ĤΔ��)aG$;9�5)����_�/�V�d�K�;����u�؏yPh*�:��:xl��ok�y�l^`UT-�Hԫ$��Sy}�n�)����I�K�Rn��+G8'�Z锆�	�	���[fS�墾c$XBz�l�,�`���O)�Kd8u.G� �0I��U���@�Xx����01�b=�̆��2E�ѳ�{?}��΁�7ϧ��;Շr �WԡU8Iyo�5�

��(&�ș�U��Z�:=����2�u��O�;�v�&�.';I�6��]m�]�M��]!X�ؕ�"G�]̳ߤe�w-m"�蓗�c��ؿ�Jvo�[ﱏ�Ǩ�mB�F���!
������}o��J�,*�*g)�ʹ�_�f>�B���N����(����ؾ��_2����V��ha���i[��$��or{�x� �Ⱡ���a��hA-��m����R-
�����<N�˘�\�`K����Q<��Y�H2 �9�0OL�gPxh����K��KO��J�9��7���[��9�SP*��=#��Q>�������Iy��wo�,pw��aܼ��=��a`*zZ;�����N\��9GN�>��8f��;�^C2ߞ��_L'��G]7w�{��r/M�[���R�$�.i� UP�lX������7t�1�Ѭ�v�u�]#aRl�]1��:L0�ա��V7���#(wp6�bH�J���][!kI ���%�ED�H��݈�y��f֥칆V���w��ľe�r�Y#wa'	d��en-�s���)oq��K�J�Xa�#��L�����81���+�Yʣ�k�$���N1�� XS�s\�~�a���YfkKPa/��.���1�����H�[���م�����x��;��P�hpg��#'(�5���?ڽLp���X�_"�&����0s�D�������H�k�"U��`���΢ѩ��c�8��_�a��x�Ҏ�8��¾��������.5��(�eac�q"��X�`猿O���*o(�#��i&���Z�܉��/������ \�:��<7Ԕ��.Tz[�0�R� �YG�b�G�V�DT��'��Z2�(̕� ���{���5�`<��͑�H�A�7t�n���D�I������
��s'{���H�S$�?w�X+g+1�	�,����V�b�x�@�vg���ˊtC�W��������?	L��8��4_7��8��)M���AS���M@���<.�e-��^3�V�����;���#�}�X^�Y�����Rb�{w�6O����g�{ޮsb8Z	�xg�/(�)Y��!9Gk�����#~��`yj{�?�bg�)ha!WR��e��2��9��H�Y�.B�h�!�����͔(������`�����6�> _�%��v�k���&�����DP��߬�q�w����";�����)	�����~])����u�↿a���j���AO��Mڿ�H|=�5zoUe���oD��q� if��k,�*�3�H�N�������LJX&�������-0�^M�l����JK�^]�x����2�C��H(�]����ᵛ΢N!6�?0�u�;@o����O�XBo=�e�K����[C`�,���N ��z����da�>��QP�>���J��A����HBk����?�03/ЏD����8�W��ED�#���ĤK{��-�|,���?������J�-��%���?�o��uGӧ��Ȩ�ǯ��1�����ˆ}8B�,���ӕм�c�it�J{E����7Y/��nր\�?�SlHf�H��q��LOdy0����'�mP�a1~	&J�y�?����̜�}��be,��j=-ݼ��"��I�#�����0�. ��Uʐ�K��Mz��:9Zb�N��8'Y�܁/R��G��+?a�D�����K���{�*e�`�<!�&M����iL=U=�*��ՂGr�q[�]�G(D��f;���4t����*e�*��;q揁D%	��C��uYv���V�l���Kd�����z6��k�h<�α���qE)�Z_��q徙h+$ڊ�u��
��]<�� ;!��"1� �����6��P��ɞ�/H}8�w�2��F�y���fvܧ[�9f.��(NT�|�j��~F!�B;�s���r�'�g�O(�֓��jz�����k�to5�=9t��i��vN\6I{{��6��i+���Oe�����9�ӽ�h��J�#�n��U=���&��:ty��n��.�<�{�}�b�r �MC��&�����6ZCa��{����:b�����0�T/��1�l�¦����)g�]Xē_"�J~!)��v�I���No��˯n���ΰ'������OEM�� j�ї�s(��v�����j��J��*�u|R��1ڟB']����}:���%�}���3J�u:y^�0�J}��$I�����`�!U�P�d�"�t�*�h�A�2X
	��C�\��ڡ�\�=�����Z�ҡ�q�mn9�����urňr&Yp��H�wGO���&6{�k�˔����.���5�L	��Ij�6���Gm��c�*J�o;���֛?:��}��c��ݞgs㶷�݇}!����N���3����#����������X$ϣ�����K��]�湺�ߞLѿ����|ƹ���%�b�������%I;(��
��\�u����X-��e]��%Ǹ��F�⛉o6�|�}l c^m���h�rT9�V�K���a�m���4Ց�,�oeEW�3o�gc���J27߹PW|ډ��ߣ]�;lNp�v��Hie�Fy?l-�Q��� ����	����mvչr3>�a�����2��`5�3�,U��1w}W�]+�RT�_5W'��W�����$�� ��Zh��l�v����S�|me�D:|S�)�kX܀l�h���VKƦ\�7���w�l�:6�X��Ab?�ʤ8����-��^BD�.Dv���O��J9v�"�"!4�#�jU�Dtv�V[������l
܎�J�u��|q���HW�ƅר�y��֜���q��t�9k�`�F�o�5 �$n��ر:SA�m|����\����A��ݙ�i��]$�8��(��27�R�2Zz_f���Q��f#���?T�J�,�m�f�~�f���#���%�e��J���������ČzmVxe�o�"{�R�K�^�p��fg���KGo5�33Kj֩��T'Q=�һ4Xj6Z�X�a���]�;���m�T��SD4���������o�3t���|��gQ-�`ib��Oɓ��i�w�!�=tT��ފ�K	 a�ۘ	\��Y&���SL��k�b��h��J5Th�7[�a>9H��*�t#��|�_4d_g5���%QM������φ�!UI
2W���D�(���Ю�{�3�t������3�%%^T����������t���'�jܪ^�y�W%h��>s@}[@"�{8h�'���V]d�S��mͥ����Z�#H��^��nG(u�� �}�9�`d��#ܾZ|7����\�!CG!����}��>F[
�Z�T�$�M�`�3����Coo�i������ѤT�~��y���P�k[�#/��� �Uz��]ҧ6��&j=�ߚ���Z��_7�B�Lc���U�7xo���ۨ�k��ӎ]V�i��w�n`�h
�kE��O�澬�k|+�I��YG"�|"'�F��,$��3Gh�:��-��Nr��cZv��q����M��C�Ʃ�˘�ʼ��=�]A�ǰ;�g��q�+RdF�sx�5�꒩��,+�eo�S�<O�+��<+����5�T�<z>�&Y��*q|Ғu���s��imq7��ZoQ0 h�GW@�JG� "r܏�V�è�ٵ#�\9�f
"j����s���a ��+�@�!K7Z�S8�����W2��yȄ�HP��-t����]��ܻxdgstnp�?w�u ��FM+2c���E2�]T�U�����wI/i��&L��yKip�!�&Q�{s,���9�'P�*�����������JaT��=t��?���0��}2r4��S7�}�T����k^�{\��Cry��堩l�H�З�F?��d���Ɩ� ��`Y�5��սgr>�1���^�����Zp�)�1�g��W��'����W���%��{�njl��-����0��v�Ê$�|m#U��UE�ػb継#��'��_Q0��4|eT\M�-� ��L���������w����0���ww�3��Z�יuz��K����9��8�y�O���v���כ��K�s��]����تh7$rP��N;�L�׃O��S���
��Ϫ\�96�}2�\v��MR��P\���ݷ�=�=�]���Jz��(
>y���.Q���.�'c�Wg�i�h�S�� �t=����-^�P:+{}����HYB�.�6�������DT-��o�|M<��`��o��̷VԻ�������OO'V��6��HU���&h��>׽'b��)AJ��938nY�<�b<��N���8�[+������Gx��놮��FWL���<�)&V>k(���mh��_/ f�����;����}2�C/;���au(5BAVs��m���ꍈ��~�I󞰹lb�5۳���'<w�g����m�If̉����3,������'�<k
h�uZ���0�����V��������]o债�;mC�-�`��� ���&PY�J���,�Ͻ8@��'����4�7����w�sl� ���g��:`�-����:�]i����7k�k. ^���G`�W��y]@`%���uLX� P ��	�4Ce��û�!类�H�f7Av� v1z*��WN���v�`+��y�* ��6�^f�,"�#h.��ǰ?WP����&�v�^����2�����͓c<���d�_I��������Q��bEKkv�*�/�<n�(s�l�e����wT�h�^T��������$�}���I2����zf�ksg:6dL�-X��;<ld�{��s����e���j��	��q���n��O�%����8��ܡ�䝈� S9z�8���ô��2� }���
*V˵"o�ыr�2��_º**�]2k���8�D�v]<�����F����+���{�U�V(�	�6����8A�A�r�]��n37�PG"�h�!�8��ݸ��y��� ["�?w��@Zթ�ʟ*�5���� ^z����g���C�t������)��G�$�e����Y�ev-]yK��H�͉�����&XkW��WՎ��`Dg$��^OW�H)3տq��=�.�K�qO��09	M��c\N��`0��TL$�K�T���\������&��r?���x9YM���44�biG�:ۦz���x�D��!~0�Q��Vo�7����`��l�+oӭ�R;���AH̳2=F��ШD;�hx���#��ۼnlM(r��ނ�
3���a�����Zn�����^���O��|��}L�h�Z5:�JJ? �-��d� �B�����ê���N���}���n��m{j(�8)}cGYP-�J:e2H?6v�T�W�G�&n�m��ya�V�@��Ǆ�$�S\0�ܹ
��<X�8?|�"�
n����NOZ�<��u��F�9�?#E�����O���"�K��`�)�%��e���@�#��~��I2eԤ:1�T����к��j��c5��֧�x��N�8)g�(^0 @�I.o��jғѴR�fx���u��QSu�~�5e�n�������e�*C������k+��P)/�9��K0�����P

�e�&x<q�7���a���O����G��Җ��#._ٿ�07v����� �ώ���gA����YU�ߧZ�K.��D�Xg6S�L��k��s8��|�N�D��C�~Q<o��9��^|C�G-��UʆW��m��J�Qsɱ�¥�~�m������+{8�����0s��[^g�I2W�e��<kFv�L�ڒ��5�n�^�*�.�P]���������/��<�_�{�C��;��U{n�h�?˒�dn��R	s< ����8:^�C��Y�h�7�=$���Ӂ���	�ڰ$���:�-}�jJ�c2��^Z��)�V�4�C�\g9��79�]�=��q�|��������։0��S��䩮	��J|,t����8�J:��A���aD+vvZӝ��kH���_;��ӟ%�M9
D5��嗑jQnk�퓄5�2��I�.	�Eok�,]�C�Z�v��l�����( ��<���kBA�/��91<]����[ѩʌ��+(C���N'�&��%�%x����Jxn����3jp8>�4Oے+L����ߏA6�:U�%�SKwT�ב�M�>w�,@����b[
�&<�s�!W�����Q���M����j��g�g'r�@Y$��ď���[@��8�<W��W��ȝ�1i>�V��>�Z��\{�98�,νƹ[n�yd��HS�����4����GK��R�mR���]�=�<9��a���.'|kD*�>��)D2��f=����B$#�х���Ӗؐ�L���ׯ�Pԙ/�ȩ10��6W��Z��vC�0<�UX��x6z�C��h�JYf�\��/O��z�F���F���yĈY��"��'H���H������N���C3}��@��ibn�.����*]�MX	P���~�ʉ�kj�R��z��E��A �Y:>>r�ɉh~���w�{�a����?*hO��/��8�w�`>�����z
#�ԝ�R]2je\/Si�KA0h[3��T�� �W��k�|���FG��a�����zS M�1���zJQ�+��̹"�z�%��M��0>3�\a�MY�����<���o^Ǒ^�gV/B�.h�s�=��<U��f|� y�0)�0�&��L���G32���RR«��Us������D�FL<���M�б�h�w0A-ҵ�[u�
gp�ļE��A�K�,dn2�C����Ne�j�5jG/H�T��Ԓ�r~��^� �|&�&���T��L����X-�\*��Z$q�iEMq�]q~R�N2�b���Fv$ _&�C�C�Tcy~�6�Ή�� T��� �X-�l��n�^��d��b������&�bg���GF��ݹ;t��	޾�xn��������`�_1���?"�\ؤv��dk��F��Ѧ�t���)�ł��yu�?�`̢����7k��Z�ň2"�~ʭ��j�h��z�_�]B,%�[���+6I��LK{��^vi�Z�)cvX�FP3��ֱ�=ଜ(k�l�g�:�L�h�i�ވ�	ʯ1���e�����]��4v����ᩩ%>.�!��܊
�z�����xL�o-C�.w�����~�����yR�T�݈ݏ����j�2[y��"��XU�Iܰh���ǰ��3͎�E���	��nL�g�4�+���y�6f����;���"好��)�|�~٩]0�ϸ��d�F�)6;�Y��*v�ഹ檧�c�y����}�cj{�}���(�g3�O�������+(+._�&��kfzگ��(��f�)�@-R���KLc�8��ߓ�w�6�}�LaR� �-+CEi���D���ͺj����W�Ga�5A�n`'g����"Ŋ�����V�W�Jr.R�B`H�|`*����涔ک�) �$g2��c*�?�H�kYY3��h,$�FP'N^K+2��4����z�Z�� ���Mo���f-�6\W� ��"��َ�X�Q�s]
p�3�� ۸ ���os;�np����Z��4��Y��'M��9�&Jjmz{�ʺ"R��>�'Y߬^*�����pK_.��+�fk�#S+�tlZ�̧SsվSb�2�{�ea������^��\���c}�c�@���Ӽ0,�S|, Oy~~��f��ֶ��}{{��w2薻�nNJqt�.�B�q����X+�E��%���9��y�6^)���y�D�6����Ԏ?^���k��	pƩ�s�����?��[��Nb�wRk�1��)��4ݻ;������M+�x
����_�UOu��@Ax�4߿M)M	%v�ޫ�qo%~�ݐ��s5�}�1���T�%���f�< pG�[P�ioo/���ܻ[�Ɔ����I�g����f-�t�9k�7	�n�k�^)5��F�fc;��!��u��1�Ic�//=��Sl���>Z�u�
�O�Y0-�p�=��Ɇ�#KZ� I�$m_��{��Q�cK(�m�!jwk-8���0�C��K�М�#����_5��7�a�7z��7>���8�l
،Z�Ch��M]&o�Уʶ�0��e:=rI���@mgp�i!�pE ����~��]`e�.Ƒ�EEM��r�D���*-mj6ȃ��o����,�ʡ������e>�j�e���jl������ԝ��*U6��&�)��Ө�d'���kb��Y�"p� �N���/,=)TXn����h��
ܼ*�ɝ���_i�Ͼ�f_vs ^�B1oL�C#����������4sED�<�m��N;
�p�l��ʳ%D�s/]���L�DJrIccrK����nIj���)&	^�E<$k�&a��J2,���p��]w�G�����	�D?N��m<��'cͷJ޲�<5�c�^�
a=��W��S�2/�oT�<|n	��x"J�i�n���Т�&fXG��P�}��5J=�2����h�vZ�0`"�gf�.-�a��	���}wW�~��������Q͊�+)�8����՞v7n��np�^|ķ#q����M ��%H���W� h� �9��ED�����R���W=)��>v�of �Q�w��s�umN�t��
S�r4�*#H3���Ԕ6.���J	���z�
sx���^�b��ܞ�d�Ew���]�����]]|+�$ҙP�p�NB�,��&ˣX��Ʋ���x�� c����肬��M/[����bfn.���S�<X�/�H��΃�T'�v�y���2�ۅ��c����t��#���7��w4���lx����T�ũ�28��;~��Z�E*IXU��Xy?�`��yP�����S`#�%��FK�hy��Z("ӽ�kvv��
�v�������
iX%="�|����5����z��g��/�M�K �e�#�"��Kc �B�x��S�e�gl���o�@Al�L�6{DO��]CH~£[��@���oz)J���m-�a���xT���*����T$'��d�e��4<_�F�m\V�K� �`:_<�Y��8ܘT�� �����|�r�f���i��$d�$[N�O#��7n:
���Q#�`t�s�xJ�	|��&�eX)�T�?3�dS�pk��8T�?�i�7����#�L>� 
�'�M�����Tr㲭�#�T�i�,l��Cȥ����-��]��:J�zU5��=q��/Z8�'].���ץRE�~������aꗙ!Pkrr3h�G�뿎�Lɖ(T���#�{Dj�w9����I�`�e+?x�u2s>;��F-Z�{�:��AʆStn���UUM�5N��%ieԹ�T�.�(��mGس�t?��>a2��t�1��������ɧ���	�ث0*�-�O�E��Hb���Ɖ$��eC`�]�H0w�$�Fܹ�1���ʼt��sФ������@����̜�=إ���57wn�>4rc�����o��}����w�J�1�Y���Pm���mZ�U��y�QW�ԃ���TN0�������N�� X�a�� �䪤x�q���⫹�~��1�ېu�7n�I�^�%���jW�d����dG2���M��W��zx�9�~�ajJ���B12�n)l#���dË�N(
��_�'b�T+	� s�:C�ҁ9�{�`��J��TN�Q��m�jc��Ρ2�NWε���h�����(�f�}N����Wp��⦷�"�m�km
|XÆq�M�,{.
�ɉ����`u�-��Tn���N1,%%�˚߲��H�]Ȗ��n W���v�*���K|�RӪ�y���ü`&?��-�2����䜁��i� I����'ѶKq�p�1��7a�j����I]ɪ��{����������o�ԞW��������챊��e ���=��V�{Gg�r�\t���a)/c3��_Z��4ҩ	]�|QL�v�T#�:*��W�kL��D� ���v�C`��c��ܧZQ����C(�r[������Zn�:I�+�t3�"Fׇ��a����B�L��6�F�5j�1�ŝ��@�d���ؔ�c�Mg	���s�ϑ�v_��H˒�ڌ~�
�Yq$$ڿ��^XXȶ~,�&��j98�d�m��&�hqh7Y��􍊑Og�B�1�E��5��f[􎢼!�u|:m��Un3��h�B���E���\�}�@��AѾײ��訠/p�5ŧ]۫'0@	����$��@
D���<�nfs~>�D��\���N�3��<��"	rXd��2��_a*�ws3��Ύ��ŀF,���͆&��s§I� q�OP��7 F��ݘ�;����7(�]+Jc�_Ó��u{�$���j�b�x�s�[:_��?m�UV�T�I��v�*��Q��2���<��ԇ����J
�4(�~R!�<Q�{�T�O�����b>�����;(u�v�O��f<������Z+b�3-\�:N�O"BD�c:D�ْ�;���:�G����{�=�j����=�7)7���::D���v�������Z(��:�xo 茏iY�՗T��9ǉ���T��ja�����l�TLM��V�sN(��장�������G��Ѓ�J8��l�NC�#$�V�&�N�_��Bͩ��>�ñ'�c� 9`x+M�pH3��)�m���a>��ѩV��#��c��d�}M����&��D�N��N��[���)?S�~�%��N%���i('/f�X9��3�H�\I�݄��K�\��{�[w�Ȁ�LY~gZ��o�
����!P��H�`��[���^��{\�iA���V�IM�n���Wv{H䓷��3��`��3$���i�υQ/uZ�X"'�S�(}�@��F/�L��Q��՛���8? -E�ZDx�^��>nԄ���>I�o�~�t���4�u{®x�΀9m M��5���܈̓�[�J���nnk�>{!�Õ���M��'7����ux�NW�7UF�绐���{��**�����k�b�B���jV>~�;����A*��T[���3>��#�G�B,�v����l�+",�p������x�PiGA��8l��N�߰�jW-�՞2�V�r�mz���RQ~"�AR�<�^i؏��\�Q"�,O0���%at�)�hY�9��y��p����.9�D�Zh�ځ�0��g+����Ř�u,e�<�!b﫥m�2�7�o���q]��#���1��i��b�mu�w���3�m��Ә���?��1�� )t�D�g-O<�|��2��B�'�	m��k�O���@H*�#�mW{�NB��0����Tڻ��ר=�$�}|����r����Y� ��\�������΁�\��l��5�ȼp_�2(t�J;xK\��a���#}7`��Q�%S�X��.���.i�w�H*�\����A{�zaF��d���-��T������5-��~� T�s�n�]v����%�V|���,_7+����ݣ�g�����$V�%���J4B �"v	�᝺�i���� ��ĵ�j3���^KIh���߁�|���W�S�&h#nkL�:��[����,�`��>w�>�R<�5jx)J!b`a��v�PiR�2]��r����)c^}��SE(C���_/4׉�w��M���#��[_�������¼�1�랟j��f��)
���y��T�8��e�T>�]��4O�r)��Т_Q<���"��4L�����)^b�L{-I)Chӯx2St��>EqC����	v-�g�+u����'���ot�������	r�s���+Z<i�iL|�PF�0ӵ.�i��P�y������C�B��B ��"/�Ы�3���Q���o��쩌"��Mf�?��2������I*��
�;�1�6D�[iسĪ/��J$��6\���&�ی�n��x<�R��ʭ��l��˳zװ��IY�`�5QE�kY*=<��.�V��$o0�1�x3'���g�.O'1WT��b�c�ZQZ]����|��'%4����� �jv�c�B�'�ُ*��� f]U�.|C���H�]�E5��@�[;u��Q�c4D�Â��qpTo���L�*̙���o�M�ۭ��aߟK��2���z�d�V�Q���$�9l��?���
0����,y>�G8��Ovs����e�Z��9������yv�X1���bQC� ]g����Y+V����ʃg��/s'�?w�)a[�VT�h��x�$,�t�t���?�Bf��6��l�jp�����F�k�:��M+��l��g�Y�?�Hq1�9x���6������&Ҿkh�����dP�������孍�W�,_�I��6�p�<��p�|aa��~���S�]���o��y��7��-q�(�rZ��-�>�M��!�\�� ��RJ��V�VZ�����d��?��:�$r!����T<,��5Ȭ����12�K-!HǭK��-��lݎ_}�׋8����0ִ��.�b��c��H=s�l�J��-|��<��t;�D��#_B�s�Ҥ��QrW�� �ɐ�K��ܮg�a�ىɯPת;Ͽ+����Az{Y��j�&���9K63��NC��jߌ���V�1��u
�Z<��F�rU��0�)��z�i�"O�>[�cǥ��g�C}׉�Xa�tvŅb��WF����o9��S����r`{�~�)#M'�-��8�"����^�i�YfI��7�9Kσ�AUΝ�&�ǋ`�z���(o7 R��<'�LQF�bb���+�ꋪ�����jG���)��[?p��֪�j	잴Tַ�9E[�kŇ�?����N|c/�����>���Ĕ��0���L9d�w���x]���D�գ��ȳ��WxT��n�a��}�y����M*,m�moT"t�����pu�u��u=��Ծ���-�e��oI"��o+.c{��d�|v�
�0c+�%�v�Y�jIZ��}�i�M\ߴEܱ�;r1��K�]'� ��q�c.�u����y�X�;6�f���yLR>��ഋEKo�(��G����UJ?�H�E�ſ_�q ^�f�]zŋL�)p=�C��嫻�=���!"!b����m�>��1Ҋ��]i
�X��r�c��˓�yA�jS��'�U�Z
��Y*!V��=���� ٨���.~/�k6�̰G�D�}�zR�� �:CU%�@n����&�C�f�K��HA�_��p�e.E	��6S��!���̸۝��O|w
�@��T�,ǡ}��r�&L$�<����؅g
��:�{ťsR�;�ܦ��o|�w��Ԕ����
&GS'H�-�Wڇ��&o~�8I۫��1�O
�*6�KG�,���m5�����K��as��Ջ�;J3��)�r;���Ʃ&�]R|���4J�TE ��i�'�i�M
�M��$�@�"����NO��(�m�����42	o�X�L]�i���v�{�\$�O6��lb�^��#"�y�e<�}Qx���+�Z��^|u�4|�$�{��S'�����@	��	yq�u��B�a=,�X1P�St�f�#����qy�%�_�w_�7 $x8X�x]���r$���X��j���S���UU�Hi�jA�RJ�X�U+�H��po�^L��^2=��<���WN�e�t�
κ�O�n�1V��6��G��T>(J�t���3ݰ_m��)��eΛ��8&5T��A{�ޢy�A���?�\���9�2�>�T�Y�v�0^������@���5��ܭS��ٗ�F��X�j������Ƴ����W�ݟ*�|:#���?������'�A,Q�uL�b�J<	�|zSRM#$���8�}a��qhޭER\:'�L��B���`6I���f ��I��zZ�9O�^�<���N)[���ק �C%���o�8B��$	�q���|����Y��b �f67�V�P��"��7�<�	X�@�Z(ڄ��)��#�^�W���`'��O.l���1��Q���� ��������t0�&�Zk��b s��"3����[�����̎�u'��$4�_�Qt��Ư���,u�M�9b�ؾb�DxH�t��6��1���{���2�-��DB1k)��H���r�`\��*�@�ꜫǝ�-"y����I5
d�I4X-F=Z,^��x���:�R���Ƀ��ޥg�0_Ec�;@�u2sn��Hb;z��Pʾ4_dښb7D��8	E��E&M_^��p�����-lu���Y�;��H"ؠQ1T�J3LQ6D� �Tzx�lu���U�Ev�����٣��\ӿ-�M��X�	�Z�]P��x���{�G$�y SL���w�[�_*|����~��Ao;cS�>�X��p߼�/�_���C�Zߎ��cV�Oze����n���X&`}?��ڻ''��k9�$�0W(���C�/K�h$2�t�b賃��imS�P�b�������$H9��#h�o&���)��^{��+��&����ߝ^@z��1-v�8�[U:��*Jz�Y�����ThL��Q��)��c����f��k@5�pZ� 2��T���{=䢯�s��?Ɏ���i_���HBB�`h��0E��R(>�-�phI�6�&W�siԶ|-�l:I#mfUȈ�:@�.�;�MH&���s@�x�����C�҆���Μ\��a�Y�U�Um]�I��<���X���W%�1�FC%zM�"H����s�p�Α�y�j�7�����W�ݗ�E�r�1��/l���*L�Vc����w��K���s�x鯗��L��]_�"{=������[����w��E�o[(eͅ��Ć��9�.Sq���ÜB$�:��J��p�v}�[JT�P8#�b8��M��p. �p�y��]�|�y�w����B�n҆yg�+ݓ��'�"�IGߏ��&V9H\M򹛻Mw>𫩁a����k��B�i��M'� Ҕ� f��ix������KjL;�nN�;��J~;�>����m�]�-�aX� t֏f�©�85�_���-V����������Y��bi�/�TC��Z���N)k~|�e����79A��n�]1�4���:j`�!Uw�����tv�}�b�{a�ngi+�c0����P���Z���1Ŋ�iS�7o���/�v��l����vS��*^V��ΦYv@���6�:�16!�I	���j��O_VȕWܞ�WԜ��3��I*�1� YG�%�@��蒘���N�qɞ�)s� }i\H��bF�x=�1�6"�H/*Ͳ�?����xP���p�SI=��HSo<�7�-�p!m�r1K�<n�v�$bEw<�Y�\��g	L�v^��YsfA�q�BZ�D>�:�CƩ2v25�%�^��LD=�h�g��O�c����u�m�k	�*�t�����)'O�Kmk�q�T)vQ�{FQ� ]�M��&!fI5��zS �WxxD�[����r0�ZlQ3q���j�B�w�o8$u�\�&6Z�b_�&�!I�������9S�큣Q��`>h/s�.�j���0����.���E2h_VfaH����f1m��'[�W���������,��P s�"B�_�1�J2F}���x9���M��1��9�)����@LL��m�n�H�.K�LAѣԖ�6����mC����2j��UE	�����a��!U���<1���er�������h�)euZ�=r�M3��|��N�m���E`آ�A�k�nL�Q3�_g��Q5���'��Q�2N��
Ҷ-�1�����v�����]5�P/�xq��@���:��79�"#銡"MrSզ\-ϳF>���__L��h	B�7ۃ�2ѓT3�*}��RG�%Y�4YU��C����t��~@&fUs�
D2�6�:f.;���G���=ݓ�2��`�Qo������D�������;��a�ZƁ��F�_#4_��!E������_o*q����zr6�}g����"5��"	\�|-�P`[z��ڲ	v>�%*�+�T��^STM�NF�#�K.�=mӲ�T{��3&ҳۨϗ�������f�z]n~]�j��pd\� i$��%{�!�C��%˨�Y��U�<z����Y�0d����ʒ&�z0�eq�ǿ2覨�vW� ��Ic��H|<��W.�|�%�b	��^I,0�D��d��&�{��k3#}(!�:Ց��:��A�Ƃ���ͤ�'AO�t���B�/�ұ%��+���uqjO�¢��Q7vф`�Y��"a]�RP�Gn^��"��l�+�WsY2�#M��m���``�J.Og��w_y�̷��q��i��[��M��!n�1�x]��L�����c�k?���M��A���p�#�Sd�H��Mڏ�C+�jV ��D��i�P�U��X����]u�G-����j1�r=Z_��R��}���$`3�B2��g��KjNנ/�0FKn��;�m۫�yGNfx�m �����}b��0�i��D(ڙ ��;"���ץ�=כyaG�',E�I�)�`K���z%�7I�]<���'K��/kg�?�TК��f�I�1�M$K��6�w�h7�&�.a�#�)�tX�e�쫽I!���ǜ����>�-0��Xb��J��Ч��ԉ:+?Uט����ge�C���N��g����:$7rS���e���ʹR����o�V[������ l�S�r�&��=��d�/�nu������/O;-C����S�D�˗\h��[�����QNT���Ά����$sC�DsQ4J��O���~>�[�_�S��r�rby��z|�免D~�Z+M֧�?�%��G��^1xv��A�z-�\A���2�?��{XA��lp4��2��/�#�r$⢺$|����M��N�D�������N �D�>g��� L|���������h�!LҸ��JFw3��/��(fVJ9[�����L�t4y��9և���k���G��}�iζbUg��T8%��e$.i���<�s��-�oLX6@0�,!� ׉���$�!�U�	�t�����Ӭc=Y��<n�w�D�̟��W
r�pQ���!��?1���ew̌�z��!g�j(&�m;�O��bF��scc�*�F��k����gM���9 a�B`����m�]��`$)~�A���P����-�b���l.��UF�i/IK�x�I�2I���r�[&�l%���(1��P,���4�# �h��~ޫY�Z������~B����RĹ���%X����y�R��Y�}��a�M�7cn&�gةP=ě'���_ %���8'����WO�����sk�W�M#��(K&�s���O�X��L$��0�#_D����5��A��:�����]��c�����8��& g����zAh���1��r:C6�L���F5�jx����\����̷S��	�J�	����5����r�7�~�K>j��|����$�A�W�w��[m��COT{�E��Bg�%�V�;͔�>�a-���X�1k1�K��S���d�)��]����<J��`�FV`f�pv��p���e���T�ePH�+�w��K'��l_�뉃�Z�� i�} ���I�����4I�$d��>e�ڂyi������&<`0|�H�l?�	ΏBYP�[�JЖ�o�V�Z�O�u����A��?+�i^���}���$JƱc4]�U�b����K����%�[��)W�x���l�zf.ۙ�x���X�\~PP&������AY�r~�d��	���E��v(��P�ߢ� S9!�T#�4�ЮC=��<��C�Cw����-��8ķ��JCF��ɸb��,��`ұm�ڥ���|*�����nT��_�uj0�$+���ޒէ������&����EV�-��*ڌ:tV��m �� �$�i�^̅?'�^�Ǡ��cHt�{5�S,>�9���.	S�߰��?���%�t�U:W�o]�F������Rt�� Ab���.�ԯG6�'Tn%���������D[���|�Gc�n�pvU�$��Ĳ���2��������������8��b�������^)Σ�u��.��S��	g=���U+T�(�l��=��>#��֭�%#&:�kwL����=ȳ<��M�[��:��|2�LM�h$]=M��e�2e���q���n�FCn��p�%x6+��%�?����������N��q����I
���:�qK���ɚC�u��u+f���eQ��ņ���� xz��q��|l�C4���hhU(������f�xM�k����3˲�~���VV&BRĻ����@������h��'ǕNN�n�.蠡J;v�/p�Զ�/U>۴�������n�s�j��m[�o���v�ma�7���t�t@�����	�-{�n�59��h�OC*�'���[��b5���p?^x5��Ҿ �� <D��f�7�}�!-F�AnS�^hnc�E7n�]'O�5:�a{��Ģ��C��B�yd�W)���*>�1{�֒�6"�Y5W2���7��.	v��ᬰ~��9tqr#3��o*��}�h��J����9wV�5QMŚ����r �<k9���lP�:�+㭣s(ʑ�jP��'��m�D#����n/e!\,�8on��Ӿ������vź(�BY�'��!�?nj�GI�Dُ�No.���0=m�$�����_C��)��9��ߢ�0:fX��ع�1���=|��B���0^=�9��ﺡ W\`]��d�R�_�׹��.2��vB���	�
v�8)��P�".l�rߪAH�v�M�a����~\LB�
f�!�le50����q�g�A�+�gv���<������ܽ^�tÁ&�}E/�f6��6�q���,D�l~��֫��j�K���~l��n������w�����wPON����7$��H�"�Q J�|��U��L\[o���1/�/%�Y���#%W�4E&��r� r�C,����wq�`�_-����{�HٻV��zI�K'��\�OO���ߎ�%|ܬ���y�;�64"����U�u���d��DJp��($i�Ϣ����6S窧P�;E=
����>��������O�"
���>AA��]��436����?��2V��G�+x��v�~��WV�d�oV�|�9李Rkӵb�p�Ϛ��6������ᄘ��8۸'q�=����p���Cx8(e9)�ѩ1s��~��v�U�I��7��1��m�.�����`�\?��-��y(�+�7��Ѷߌ���cˁv��!���Taˉv����y�s&��b�	���
ɛ���w�#������bA��ۭ)��r�٧��{g�i�eS��_����|���G~=�}��iv�v2�>��x�1��Uy��o� -��nP,����0��8��X�W��S���z��,'�MG��=�����߾:o�o��?'Z=�-��,�1��y���mn�\�-WK�����<�Ǌ?x��޿O�M�B�b-��L�X#ԏ�~��dB������'���V��j�r$

��e6`#��t�V���ԾlW�]��I%�d_N|&g�Z�=t����l��ԉ��hp {t,}���(3zXw9��Q�Ϋ���>L�r�F�ɵ
�ß�RB�hr��Uto����3j�����AI���xVXPa�Ngwe���?��~/}��Ұ���g�!~`7a�D�|ᰩ?Uހ�bȞ�?�:��G*Fj"Ӫ�bw���,^�P����j�u&�v�)�@���#���ٽ�eI$�	��/|�.�z�9�h-��5��3rL�֔���g#������\����8:'܅,ө
���~.A�
��h��b�k�9����U{�tvo,��j�ؚrq5ǩI��;v�aDؗ^��Qw���z�����|�O��y�:LS�"7�)'�ԵԨ^>���B��წ{�נA����kK+���ީl*�[�Z2Mҽ�=��ӭɫ��Rh�d\�S>z��S�ff|���1d���V	y��rJ�>�����x�s_�Ʃ�����qz�m+�l�O��¿.��ON���4�K��b�v�ˑ�n���K�R�B�?S���������PX7������n3��sW�`]�dX����ӱ`h�R<j�`�O�����L���à��c.��y�q�g���&���H`c�}?X��%�_8J�o�;�0�@!�!��Z:��������I� �3�a>��+�O��W���+4��89wG�I�)*5�N�$]���� ���?�|S8cރ����8d/��j��9c	�yV/x(������^�`)���d6�bz�E�o�r�j�2���_��Q:k%\�����)ե��3�	��lv�~�A5�%���nH��v�V�����"mǵ&�&7�޹}j���e=LO0��͜��a\���/�p�LI��f^i�!�ഝ�R�pJ��
A�#�ֳv�n^��o4������y���=��.��"LM�G��G���>������H�:���i;}y��q���v��;�g�4�f�)���r�T��,�^��6˫$|\נ��l�q�#��ئWcP9���O��V3��z���Ǟ
m��wJ�,#��^2dHR!���0Y���&\�p�F�l��VW1�X%���4��=}���������3�s�������6�L$��M�{	7��<g��Y��c}���Z*�*����N����#-e�����n�Ǖ���Q����Z.Ps�\l@����'Xs����Z℟l.��� Q<���L��64�8H�q�n��~6��rS����Q1(���P��I�鯌f9R���m�yU���'ʒ�^�:��<��}�p��*�@��UF���_ ��O����|�:$�`����Θ�� �(\�Uw�9���AeMv��j�g~��)�
#v�S`)&�x�-`^�j�՞�h�,�d��Ԥ#�U2��Z7v}Qǅ>E��̷؞�X�V���i���WrH
^�#]"��8x@��������}2"L'�+m�%͊*�^d�H���r5ù�6�骜��5H�¿..e��7���hq�c�\����.�w�t��(2�k^Ť�/d;���DN�֊��"�hn��v?��׶�|�:m��:�f��9t��M�~(ƃ#��'��1!�b��7�E�l]��x������^��	�/z�i��,t���!c��y
|�'9��!���z{" m[Kc�{47�ɸ�I��U��~�B^�Y����I�~�\�)v�@]e�J�ꮃT<9U��X7B���MQ�ڙ9�N21p���/��7@p���4�u��JN�h��1|�~�ԪX�DO��x�N�A�T���l�-s~-�5�sH��T��\TќY${q��9E���E����#4�b)�P��N]KnIٮ��X�^�&��@k����g��ly�q��KYaHN}�}*$�Q�n����G�n�\u�`f)�K?�\�?:7��w�=����G3��KH�~�O�*�S�;��r���c@x��)J�jl���Jߡ������Н.Д��X�:�~�r`Zp��f�/��$D+��������CZ\��w��9Fr���ԽKش�?���KA��jq�RuFn��
-��]yn����'-3 i$����X�-$����e,,�Td��^�Ὧ�բg�2�K��`;�Zb�9��S����������YB�������$Q79wi[�^$��5��4�\�1+*���?b?��)E,ߥ%�S(��_bV��|�B[6�h�\���;�@;�ތSk/(Z���� Pݳc	$�n�T��+��A���N�s�MmKk��j,���F���A3�V悂����y]�7����g늦��Lv�ߚ��	��̍ԩ�@��\C����6x^.�m���b]:b-;|��Wb֪#Az��0P4����֫�vUp%6�y��Ҫo�d��Z����Ό񠳕A{���{ğmMֲًp�> *fs���]�?��ȓXC{=ҍO���ډ5�W/�\�-.���B�wڻt�����K-l���A|]]�1�R�4�Qf�`�����^�k�R;'�b�/Qg��B��P�y9}Ռ�U�8|��ƒ��!O���XN�mo:Z }ܶ�'��Xùhe=�]9���v��!��G�*Q~�/?1{��d5��^ߊ~-q.T��� ��v��^I%By�؉h��Ew���C���^��`�[��.;��
���Η"��2G�#�3w�����uK�� s6۱w�u��t{v߽�_Xɜw�����۫2�����tP"<]��/V7�� �����n`n)>�0Ƨ\�Zoq���G6{6P�Uc��0�H\u٩�+���6�p4BḠ���q����PG�����o}3���*#Hsߣ��ӖG�s~�E3^=q~�k�Kz�����0�ҘC[��ra��� rs^��-�H�o,c]�U�����Ƙn`�| Q 51�[��{H����Ko����
w���Z�+#[RX�C����1��uJ�;���Su����c;�^ 3�������8;�?\�{��\���δ�����Jf���eu���n�.QuG��D޶��˖��3®���a�{��ԾtL��J����
���z�_¯R���ӽqb����m��@�'�[��� j�_uE����-��B���l��;�5a1�$p���`ݻ��ȧ�dX
�4&g���_k������ظ3�z�d��w���j'd�"S8��a�f����Va��c֍R��������L�&��?�^�A��Q����u�}�p��-|�8fJ��?�<�̛�))"� ���P����v(í�zF1��v����h�w��j�{F�>�H<{odX0�*�����L�~zb�04�R��B�xs���2+~�C��ٸ�ٸڇF��\��'8�E�o���Gw���ץ#�L�bv���<���/�u&�\���B//��{#��Wk��N��U�H��Mb��ɨA����G~�/�4�!�U�W��3��Rz��̺訩3\;�t.����r�ry�t�N��!2WC��]�l�Z��a�n�jј�S n��Q��ݺ��~V�Uhs�Ĕ��F�I3v��X�~�nVu�(�_ F셄�I�������B�j�k��wgM�����:>o��W����'DdU��M�����S1jw�3�9-1;-�Mf{��8�v�cԪ�M�^�_��\Dg��D�a�!��+Dz! �c�L�Ѧ��Gmv�ᇠ�|��>+x�U	�?z���S�//ص\�׫��FIfS{=E�_�n���Xb�GG�N4�rka��uU>iE/[���A��9�z=!|d�8F�xd�n��9�9l���ۧ��]b/VPs�iӈ-!�ᱵ��kH���a�Β��.x�����
�N�x28j�VF�ב.ro�@7��������S�ը9�4F�?I<�zm�=�"ボ�g�H�5hN�d���m%�ݫ�p�	o<��sn���D1|O)�<��e.�K�$��o��/��C%��!M�	,��1����-��Y˹>�V����Ok�NO�E�4�䲂���(>�I,��ʧ$����E�_o~}��d_HT-��l$y�,:�;C#s��ҳM="�-1Fι'�ᷬ7�LW�!O����~���gƩ���l<39!��	�ڗ�Z�)�j_X���0&��z�,7��-i|>�ܓ`�ZL�ո�!�����5j��:+ZΘJYp]V��o�Jyx��1'�.f/�]�?|��Sy=r�K��-l����xZ䖭�v�^d�+(]]/m��tQW?P��;
��K�|��r��"=��GIp����q�W�'O]8.kX�.&���ewt�6�*$0Ю�w# � -���̾�� �k������<�� )�W�a��3�~:�3����-*ymo��:g0jz��k�4Z�g-�.Gzn[mU-i.k��Y�]n���W6Y����
	���O4~'RN�LW�� ���\�ǧ��"j��d(c��9*���PM:e��瀎y�߂C�U?�OSݳ9hA.�4��!_�1p��g�-"�܄baw���}-:s��i�Ml��E���Pʰ���~���qn�	�)���&����+y%F��ᄸW�'5bP�M�T��uyB\�����]����V��#4��9�YM�uhq�9�#8.��cȂ���&�g0?�_�*(�+[{{D�o�>�4I�\u#ĭ���SY��Gۙ��k�g�`���{P{?4�_�kq�bg~㋱���g�6���%��~ւtE���Ok��q/��9Tf�JBq�t�����τ�ѳ�,6����WjQ��.Z~�0R��r=��(F	����H�(c
��k4�幨K֣F��i��Tz S�4�__'��̂�������r�΂���(P\)��7�I23WpZ̾�_̤\�Yy�3�Δ�t���ف�+�.��w�b�H���t�q��7f�
�|��:5Q�%�y�z^<��`vd�%��� ���Jf��h�w��H_���>͓i�� ��e���8$�J?�f���H����R]ge�J�v�D��r�ύ`2��=Y���'\1���1 ,J��d�e�(VDTK���7�#��N�������)�[R/�nNh�sz�&k���w��j������A����>7<������a����*���\ˍ��o00&�)���_<u`��	�B��GO�pvOP/���JLgA!�p65����q��������%o+�>�{j�������PK   ¬eX��xV  �     jsons/user_defined.json���n�6�_%�U�����"�F����E��(*�H�lwy��	�-M�j�l��G���<g����.����_*_7���Y���wM���!��dw(������?���0��ꆳ�8\l��G늽���'�-ڽ�[����ۇ���ew�#n�J���?����º�#e��"
*��h�
��S�}3s�s}�ݟv����q����'K�+�0ZST%��B0&U����y����IƂ�H�dM�7�U�,�U^}��X��_;<쉿���/�p�b(m�e��Y{x�7��x��6��ɜK�{���(ϭ�ƞ�8���6�T�Z�{�ᐗa@�k��f3�ʸ���(g<W�
3�s��u]���b�)J?L�x���ίO��)������u������X ��������� � �V(��s%���1�(��d� C��,h��)%�� 0�Z6���8�AY���ţdB �,L�SQ�	���f�t\o��9(.-L �x��P҃��l�h��h��A
��S�Z���=H0bB����	��=H���a�Ϣ�P�غU���L����_Ki$H��_{7�60��3��U3FE*��w��(�X��+�
X��z(U��J>�������ع������( T�qS���� ��������7mv�~f\�FK��"�W);s=S�9�oiz� B![#r��L��x�f����Zu��#�E�1��S���H~C+�>�T%7��F�B	�>ɓˇ������oO>�kӣ%y�G}����9:��m��v�~�Ft���Nh��bN�W��]���3>�QSi��-	0W(���*+�+����}�� HY%�u,)������
P ����
���W'�_b�,���k�kex���6@��Yプ,���D�c��WQ�W��u�߳��`|��>jF��Ga��~�`|�	 d:����b��'�f���	�G�֦��&~P��c���7�	 y:`���b{N � ����P����PK
   ¬eX�n�  �                   cirkitFile.jsonPK
   �eX��D>  ?>  /               images/3d2da6db-3dc1-43d2-90bb-751371ef683b.pngPK
   �eX�C��z �� /             �K  images/a1fe0c5b-edee-4877-8adb-d45444225416.pngPK
   �eX�����"  �"  /             �� images/a890ee50-b65f-4e8d-9ddc-5b796e5840d1.pngPK
   �eX� ��! �3 /             � images/adef7304-bf01-4449-bba8-564470ca0600.pngPK
   ¬eX��xV  �               7 jsons/user_defined.jsonPK      �  t   